VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
	DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.02 ;

USEMINSPACING OBS OFF ;

CLEARANCEMEASURE MAXXY ;


PROPERTYDEFINITIONS 
END PROPERTYDEFINITIONS
LAYER ACTI

	TYPE MASTERSLICE ;
END ACTI

LAYER POLY

	TYPE MASTERSLICE ;
END POLY

LAYER CONT

	TYPE CUT ;
	SPACING 0.6  ;
	SPACING  0.6 
		SAMENET LAYER  CONT ;

END CONT

LAYER MTL1

	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
	PITCH 1.32 ;
	WIDTH 0.48 ;
	OFFSET 0 ;
	SPACING 0.52  ;
	SPACING  0.52 
		SAMENET ;

	WIREEXTENSION 0.24 ;
	MAXWIDTH 2.14748e+06 ;
	MINWIDTH 0.48 ;
	RESISTANCE RPERSQ 0.044 ;
	CAPACITANCE CPERSQDIST 2.5e-05 ;
	THICKNESS 0.5 ;
	MINIMUMDENSITY 30 ;
	MAXIMUMDENSITY 70 ;
	ANTENNAMODEL OXIDE1 ;
	ANTENNAAREARATIO 5000 ;
END MTL1

LAYER VIA1

	TYPE CUT ;
	SPACING 0.6  ;
	
END VIA1

LAYER MTL2

	TYPE ROUTING ;
	DIRECTION VERTICAL ;
	PITCH 1.44 ;
	WIDTH 0.48 ;
	OFFSET 0.72 ;
	SPACING 0.52  ;
	SPACING  0.52 
		SAMENET ;

	WIREEXTENSION 0.24 ;
	MAXWIDTH 2.14748e+06 ;
	MINWIDTH 0.48 ;
	RESISTANCE RPERSQ 0.037 ;
	CAPACITANCE CPERSQDIST 1.6e-05 ;
	THICKNESS 0.5 ;
	MINIMUMDENSITY 30 ;
	MAXIMUMDENSITY 70 ;
	ANTENNAMODEL OXIDE1 ;
	ANTENNAAREARATIO 5000 ;
END MTL2

LAYER VIA2

	TYPE CUT ;
	SPACING 0.6  ;
	
END VIA2

LAYER MTL3

	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
	PITCH 1.32 ;
	WIDTH 0.64 ;
	OFFSET 0 ;
	SPACING 0.6  ;
	SPACING  0.6 
		SAMENET ;

	WIREEXTENSION 0.32 ;
	MAXWIDTH 2.14748e+06 ;
	MINWIDTH 0.64 ;
	RESISTANCE RPERSQ 0.027 ;
	CAPACITANCE CPERSQDIST 1.1e-05 ;
	THICKNESS 0.5 ;
	MINIMUMDENSITY 30 ;
	MAXIMUMDENSITY 70 ;
	ANTENNAMODEL OXIDE1 ;
	ANTENNAAREARATIO 5000 ;
END MTL3

LAYER VIA3

	TYPE CUT ;
	SPACING 1.56  ;
	
END VIA3

LAYER MTL4

	TYPE ROUTING ;
	DIRECTION VERTICAL ;
	PITCH 3.24 ;
	WIDTH 1.44 ;
	OFFSET 0 ;
	SPACING 1.4  ;
	SPACING  1.4 
		SAMENET ;

	WIREEXTENSION 0.72 ;
	MAXWIDTH 2.14748e+06 ;
	MINWIDTH 1.44 ;
	RESISTANCE RPERSQ 0.027 ;
	CAPACITANCE CPERSQDIST 1.1e-05 ;
	THICKNESS 0.8 ;
	MINIMUMDENSITY 25 ;
	MAXIMUMDENSITY 70 ;
	ANTENNAMODEL OXIDE1 ;
	ANTENNAAREARATIO 5000 ;
END MTL4

VIARULE VIAGEN12 GENERATE 
	LAYER MTL2 ;
		ENCLOSURE 0.12 0.12 ; 
		WIDTH 0 TO 1000 ;
	LAYER MTL1 ;
		ENCLOSURE 0.12 0.12 ; 
		WIDTH 0 TO 1000 ;
	LAYER VIA1 ;
		RECT -0.2 -0.2 0.2 0.2 ;
		SPACING 1 BY 1 ;

END VIAGEN12 

VIARULE VIAGEN21 GENERATE 
	LAYER MTL1 ;
		ENCLOSURE 0.12 0.12 ; 
		WIDTH 0 TO 1000 ;
	LAYER MTL2 ;
		ENCLOSURE 0.12 0.12 ; 
		WIDTH 0 TO 1000 ;
	LAYER VIA1 ;
		RECT -0.2 -0.2 0.2 0.2 ;
		SPACING 1 BY 1 ;

END VIAGEN21 

VIARULE VIA2GEN23 GENERATE 
	LAYER MTL3 ;
		ENCLOSURE 0.2 0.2 ; 
		WIDTH 0 TO 1000 ;
	LAYER MTL2 ;
		ENCLOSURE 0.12 0.12 ; 
		WIDTH 0 TO 1000 ;
	LAYER VIA2 ;
		RECT -0.2 -0.2 0.2 0.2 ;
		SPACING 1 BY 1 ;

END VIA2GEN23 

VIARULE VIA2GEN32 GENERATE 
	LAYER MTL2 ;
		ENCLOSURE 0.12 0.12 ; 
		WIDTH 0 TO 1000 ;
	LAYER MTL3 ;
		ENCLOSURE 0.2 0.2 ; 
		WIDTH 0 TO 1000 ;
	LAYER VIA2 ;
		RECT -0.2 -0.2 0.2 0.2 ;
		SPACING 1 BY 1 ;

END VIA2GEN32 

VIARULE VIA3GEN43 GENERATE 
	LAYER MTL3 ;
		ENCLOSURE 0.32 0.32 ; 
		WIDTH 0 TO 1000 ;
	LAYER MTL4 ;
		ENCLOSURE 0.4 0.4 ; 
		WIDTH 0 TO 1000 ;
	LAYER VIA3 ;
		RECT -0.72 -0.72 0.72 0.72 ;
		SPACING 3 BY 3 ;

END VIA3GEN43 

VIARULE VIA3GEN34 GENERATE 
	LAYER MTL4 ;
		ENCLOSURE 0.4 0.4 ; 
		WIDTH 0 TO 1000 ;
	LAYER MTL3 ;
		ENCLOSURE 0.32 0.32 ; 
		WIDTH 0 TO 1000 ;
	LAYER VIA3 ;
		RECT -0.72 -0.72 0.72 0.72 ;
		SPACING 3 BY 3 ;

END VIA3GEN34 

VIA CON_MA 
	RESISTANCE 14 ;
	LAYER ACTI ;
		RECT -0.36 -0.36 0.36 0.36 ;
	LAYER CONT ;
		RECT -0.2 -0.2 0.2 0.2 ;
	LAYER MTL1 ;
		RECT -0.32 -0.32 0.32 0.32 ;

END CON_MA 

VIA CON_MM3 DEFAULT 
	RESISTANCE 8 ;
	LAYER MTL3 ;
		RECT -1.04 -1.04 1.04 1.04 ;
	LAYER VIA3 ;
		RECT -0.72 -0.72 0.72 0.72 ;
	LAYER MTL4 ;
		RECT -1.12 -1.12 1.12 1.12 ;

END CON_MM3 

VIA CON_MP 
	RESISTANCE 8 ;
	LAYER POLY ;
		RECT -0.36 -0.36 0.36 0.36 ;
	LAYER CONT ;
		RECT -0.2 -0.2 0.2 0.2 ;
	LAYER MTL1 ;
		RECT -0.32 -0.32 0.32 0.32 ;

END CON_MP 

VIA DCON_MM2_east DEFAULT 
	RESISTANCE 0.35 ;
	LAYER MTL2 ;
		RECT -0.32 -0.32 1.32 0.32 ;
	LAYER VIA2 ;
		RECT -0.2 -0.2 0.2 0.2 ;
		RECT 0.8 -0.2 1.2 0.2 ;
	LAYER MTL3 ;
		RECT -0.4 -0.4 1.4 0.4 ;

END DCON_MM2_east 

VIA DCON_MM2_north DEFAULT 
	RESISTANCE 0.35 ;
	LAYER MTL2 ;
		RECT -0.32 -0.32 0.32 1.32 ;
	LAYER VIA2 ;
		RECT -0.2 -0.2 0.2 0.2 ;
		RECT -0.2 0.8 0.2 1.2 ;
	LAYER MTL3 ;
		RECT -0.4 -0.4 0.4 1.4 ;

END DCON_MM2_north 

VIA DCON_MM2_south DEFAULT 
	RESISTANCE 0.35 ;
	LAYER MTL2 ;
		RECT -0.32 -1.32 0.32 0.32 ;
	LAYER VIA2 ;
		RECT -0.2 -1.2 0.2 -0.8 ;
		RECT -0.2 -0.2 0.2 0.2 ;
	LAYER MTL3 ;
		RECT -0.4 -1.4 0.4 0.4 ;

END DCON_MM2_south 

VIA DCON_MM2_west DEFAULT 
	RESISTANCE 0.35 ;
	LAYER MTL2 ;
		RECT -1.32 -0.32 0.32 0.32 ;
	LAYER VIA2 ;
		RECT -1.2 -0.2 -0.8 0.2 ;
		RECT -0.2 -0.2 0.2 0.2 ;
	LAYER MTL3 ;
		RECT -1.4 -0.4 0.4 0.4 ;

END DCON_MM2_west 

VIA DCON_MM_east DEFAULT 
	RESISTANCE 0.35 ;
	LAYER MTL1 ;
		RECT -0.32 -0.32 1.32 0.32 ;
	LAYER VIA1 ;
		RECT -0.2 -0.2 0.2 0.2 ;
		RECT 0.8 -0.2 1.2 0.2 ;
	LAYER MTL2 ;
		RECT -0.32 -0.32 1.32 0.32 ;

END DCON_MM_east 

VIA DCON_MM_north DEFAULT 
	RESISTANCE 0.35 ;
	LAYER MTL1 ;
		RECT -0.32 -0.32 0.32 1.32 ;
	LAYER VIA1 ;
		RECT -0.2 -0.2 0.2 0.2 ;
		RECT -0.2 0.8 0.2 1.2 ;
	LAYER MTL2 ;
		RECT -0.32 -0.32 0.32 1.32 ;

END DCON_MM_north 

VIA DCON_MM_south DEFAULT 
	RESISTANCE 0.35 ;
	LAYER MTL1 ;
		RECT -0.32 -1.32 0.32 0.32 ;
	LAYER VIA1 ;
		RECT -0.2 -1.2 0.2 -0.8 ;
		RECT -0.2 -0.2 0.2 0.2 ;
	LAYER MTL2 ;
		RECT -0.32 -1.32 0.32 0.32 ;

END DCON_MM_south 

VIA DCON_MM_west DEFAULT 
	RESISTANCE 0.35 ;
	LAYER MTL1 ;
		RECT -1.32 -0.32 0.32 0.32 ;
	LAYER VIA1 ;
		RECT -1.2 -0.2 -0.8 0.2 ;
		RECT -0.2 -0.2 0.2 0.2 ;
	LAYER MTL2 ;
		RECT -1.32 -0.32 0.32 0.32 ;

END DCON_MM_west 

VIARULE TURN1 
	LAYER MTL1 ;
		DIRECTION HORIZONTAL ;

END TURN1 

VIARULE TURN2 
	LAYER MTL2 ;
		DIRECTION HORIZONTAL ;

END TURN2 

VIARULE TURN3 
	LAYER MTL3 ;
		DIRECTION HORIZONTAL ;

END TURN3 

VIARULE TURN4 
	LAYER MTL4 ;
		DIRECTION HORIZONTAL ;

END TURN4 

SITE standard 
	CLASS CORE ;
	SYMMETRY Y ;
	SIZE 1.44 BY 13.2 ;
END standard 

SITE blocksite 
	CLASS CORE ;
	SYMMETRY X Y R90 ;
	SIZE 0.1 BY 0.1 ;
END blocksite 

SITE tp_iosite 
	CLASS CORE ;
	SYMMETRY Y ;
	SIZE 0.1 BY 400 ;
END tp_iosite 

SITE tp_cornersite 
	CLASS CORE ;
	SYMMETRY X Y R90 ;
	SIZE 400 BY 400 ;
END tp_cornersite 

SITE bp_iosite 
	CLASS CORE ;
	SYMMETRY Y ;
	SIZE 0.1 BY 190 ;
END bp_iosite 

SITE bp_cornersite 
	CLASS CORE ;
	SYMMETRY X Y R90 ;
	SIZE 190 BY 190 ;
END bp_cornersite 

MACRO VDDTIE
	CLASS CORE ;
	FOREIGN VDDTIE 0 0  ;
	ORIGIN 0 0 ;
	SIZE 2.88 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 8.92 1.12 11.22 ;

		END 

		ANTENNADIFFAREA 2.112 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 2.88 13.68 ;
			RECT 1.8 9.04 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 2.88 1.46 ;
			RECT 0.48 -0.48 1.12 2.28 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.48 3.26 2.16 3.92 ;
			RECT 1.48 3.26 2.16 4.92 ;

	END

END VDDTIE

MACRO TLATX3
	CLASS CORE ;
	FOREIGN TLATX3 0 0  ;
	ORIGIN 0 0 ;
	SIZE 24.48 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN E
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 3.96 1.04 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.907 LAYER MTL1  ;
	END E
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 2.48 7.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.907 LAYER MTL1  ;
	END SE
	PIN CK
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 7.86 9.68 8.34 ;
			RECT 9.04 3.14 9.68 8.34 ;
			RECT 8.4 3.14 9.68 3.78 ;
			RECT 7.6 7.86 8.24 8.5 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.936 LAYER MTL1  ;
	END CK
	PIN ECK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 23.44 7.44 24.08 11.22 ;
			RECT 20.64 7.44 24.08 7.92 ;
			RECT 22 3.82 22.64 7.92 ;
			RECT 20.52 3.82 22.64 4.3 ;
			RECT 20.64 7.44 21.28 11.22 ;
			RECT 20.52 1.98 21.16 4.3 ;

		END 

		ANTENNADIFFAREA 8.37 LAYER MTL1  ;
	END ECK
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 24.48 13.68 ;
			RECT 22.04 8.44 22.68 13.68 ;
			RECT 19.2 9.02 19.84 13.68 ;
			RECT 16.4 9.06 17.04 13.68 ;
			RECT 13.28 10.22 14.92 13.68 ;
			RECT 8.04 9.5 8.68 13.68 ;
			RECT 2.8 9.7 3.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 24.48 1.46 ;
			RECT 21.92 -0.48 22.56 3.26 ;
			RECT 19.08 -0.48 19.72 2.94 ;
			RECT 15.04 -0.48 15.68 2.42 ;
			RECT 8.92 -0.48 9.56 2.62 ;
			RECT 3.68 -0.48 4.32 2.34 ;
			RECT 0.4 -0.48 1.04 2.62 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 2.04 1.98 2.68 3.34 ;
			RECT 2.04 2.86 4.68 3.34 ;
			RECT 4.04 2.86 4.68 9.18 ;
			RECT 0.4 8.7 4.68 9.18 ;
			RECT 0.4 8.7 1.04 11.22 ;
			RECT 5.6 1.98 6.72 2.62 ;
			RECT 5.6 1.98 6.32 5.78 ;
			RECT 5.6 1.98 6.08 11.22 ;
			RECT 5.2 9.58 6.08 11.22 ;
			RECT 7.24 1.98 8.16 2.62 ;
			RECT 7.24 1.98 7.72 7.14 ;
			RECT 7.04 3.14 7.72 7.14 ;
			RECT 6.6 6.5 8.52 7.14 ;
			RECT 6.6 6.5 7.08 10.14 ;
			RECT 6.6 9.5 7.3 10.14 ;
			RECT 10.2 1.98 11 3.78 ;
			RECT 10.2 3.14 11.48 3.78 ;
			RECT 10.2 1.98 10.68 11.22 ;
			RECT 9.46 9.02 10.68 11.22 ;
			RECT 11.8 1.98 12.48 2.62 ;
			RECT 12 1.98 12.48 5.78 ;
			RECT 11.2 5.14 12.84 5.78 ;
			RECT 11.36 5.14 11.84 9.22 ;
			RECT 11.2 8.58 11.84 9.22 ;
			RECT 13.8 3.42 15.68 4.06 ;
			RECT 13.8 3.42 14.64 8.86 ;
			RECT 12.64 7.22 14.64 8.86 ;
			RECT 14 3.42 14.64 9.34 ;
			RECT 15.48 5.86 18.96 6.34 ;
			RECT 15.48 5.86 16.12 7.5 ;
			RECT 18.32 5.86 18.96 7.5 ;
			RECT 16.68 2.14 17.32 5.3 ;
			RECT 16.68 4.82 20.32 5.3 ;
			RECT 19.48 4.82 20.32 6.46 ;
			RECT 19.48 4.82 19.96 8.5 ;
			RECT 17.8 8.02 19.96 8.5 ;
			RECT 17.8 8.02 18.44 11.22 ;

	END

END TLATX3

MACRO TINV3
	CLASS CORE ;
	FOREIGN TINV3 0 0  ;
	ORIGIN 0 0 ;
	SIZE 18.72 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 9.48 4.96 11.12 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 8.986 LAYER MTL1  ;
	END A
	PIN EN
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 3.96 3.92 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 3.269 LAYER MTL1  ;
	END EN
	PIN O
		DIRECTION OUTPUT TRISTATE ;
		PORT 
			LAYER MTL1 ;
			RECT 16.56 7.38 17.2 10.02 ;
			RECT 10.68 7.38 17.2 7.86 ;
			RECT 13.64 7.38 14.28 10.02 ;
			RECT 11.92 2.98 12.56 7.86 ;
			RECT 10.68 7.38 11.32 10.02 ;

		END 

		ANTENNADIFFAREA 13.392 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 18.72 13.68 ;
			RECT 7.72 9.12 8.36 13.68 ;
			RECT 4.76 9.12 5.4 13.68 ;
			RECT 1.8 10.34 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 18.72 1.46 ;
			RECT 9.08 -0.48 9.72 3.44 ;
			RECT 6 -0.48 6.64 4.54 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 4.28 1.98 4.92 2.62 ;
			RECT 4.44 1.98 4.92 7.6 ;
			RECT 4.28 6.96 5.92 7.6 ;
			RECT 2.28 7.12 5.92 7.6 ;
			RECT 2.28 7.12 2.76 9.82 ;
			RECT 0.4 9.34 2.76 9.82 ;
			RECT 0.4 9.34 1.04 10.98 ;
			RECT 10.52 1.98 14.24 2.46 ;
			RECT 7.4 2.96 8.04 4.44 ;
			RECT 10.52 1.98 11.16 4.44 ;
			RECT 7.4 3.96 11.16 4.44 ;
			RECT 13.6 1.98 14.24 4.54 ;
			RECT 3.28 8.12 9.8 8.6 ;
			RECT 3.28 8.12 3.92 10.02 ;
			RECT 6.24 8.12 6.88 10.02 ;
			RECT 9.16 8.12 9.8 11.22 ;
			RECT 12.16 8.38 12.8 11.22 ;
			RECT 15.12 8.38 15.76 11.22 ;
			RECT 9.16 10.74 15.76 11.22 ;

	END

END TINV3

MACRO TINV2
	CLASS CORE ;
	FOREIGN TINV2 0 0  ;
	ORIGIN 0 0 ;
	SIZE 11.52 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 5.96 8.24 7.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 4.637 LAYER MTL1  ;
	END A
	PIN EN
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.72 4.96 5.36 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.757 LAYER MTL1  ;
	END EN
	PIN O
		DIRECTION OUTPUT TRISTATE ;
		PORT 
			LAYER MTL1 ;
			RECT 10.32 8.12 11.12 11.22 ;
			RECT 10.48 1.98 11.12 11.22 ;
			RECT 7.48 8.12 11.12 8.6 ;
			RECT 7.48 8.12 8.12 10.22 ;

		END 

		ANTENNADIFFAREA 9.008 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 11.52 13.68 ;
			RECT 4.68 9.12 5.32 13.68 ;
			RECT 1.8 10.34 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 11.52 1.46 ;
			RECT 7.8 -0.48 8.44 4.54 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 4.2 6.96 6.72 7.6 ;
			RECT 6.08 1.98 6.72 7.6 ;
			RECT 2.24 7.12 6.72 7.6 ;
			RECT 2.24 7.12 2.72 9.82 ;
			RECT 0.4 9.34 2.72 9.82 ;
			RECT 0.4 9.34 1.04 10.98 ;
			RECT 3.24 8.12 6.72 8.6 ;
			RECT 6.08 8.12 6.72 11.22 ;
			RECT 3.24 8.12 3.88 11.22 ;
			RECT 8.88 9.12 9.52 11.22 ;
			RECT 6.08 10.74 9.52 11.22 ;

	END

END TINV2

MACRO TINV
	CLASS CORE ;
	FOREIGN TINV 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 6.22 6.8 7.86 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.246 LAYER MTL1  ;
	END A
	PIN EN
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.84 4.96 2.48 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.166 LAYER MTL1  ;
	END EN
	PIN O
		DIRECTION OUTPUT TRISTATE ;
		PORT 
			LAYER MTL1 ;
			RECT 6.08 8.92 6.8 11.22 ;
			RECT 4.72 3.42 6.8 3.9 ;
			RECT 6.16 1.98 6.8 3.9 ;
			RECT 4.72 8.92 6.8 9.56 ;
			RECT 4.72 3.42 5.36 9.56 ;

		END 

		ANTENNADIFFAREA 5.635 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 2.68 10.56 4.32 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 3.76 -0.48 4.4 2.62 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 2.12 1.98 3.24 2.62 ;
			RECT 2.76 1.98 3.24 3.62 ;
			RECT 1.8 7.22 3.48 7.86 ;
			RECT 3 3.14 3.48 10.04 ;
			RECT 0.84 9.56 3.48 10.04 ;
			RECT 0.84 9.56 1.48 10.98 ;

	END

END TINV

MACRO SCHMTTE
	CLASS CORE ;
	FOREIGN SCHMTTE 0 0  ;
	ORIGIN 0 0 ;
	SIZE 15.84 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.04 4.96 5.68 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 3.182 LAYER MTL1  ;
	END A
	PIN EN
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.72 6.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.267 LAYER MTL1  ;
	END EN
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 13.4 7.98 15.44 8.46 ;
			RECT 14.8 1.98 15.44 8.46 ;
			RECT 13.4 7.98 14.04 10.62 ;

		END 

		ANTENNADIFFAREA 4.467 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 15.84 13.68 ;
			RECT 14.8 8.98 15.44 13.68 ;
			RECT 12.4 4.3 13.12 5.94 ;
			RECT 12.4 4.3 12.88 10.02 ;
			RECT 12 9.54 12.64 13.68 ;
			RECT 2.72 8.44 3.36 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 15.84 1.46 ;
			RECT 11.4 3.3 14 3.78 ;
			RECT 13.36 -0.48 14 3.78 ;
			RECT 11.08 8.26 11.88 8.9 ;
			RECT 11.4 3.3 11.88 8.9 ;
			RECT 0.48 -0.48 1.12 4.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 4.68 2.18 5.5 2.82 ;
			RECT 4.68 2.18 5.16 4.44 ;
			RECT 4.52 3.8 5.16 4.44 ;
			RECT 6.16 3.8 7.44 4.44 ;
			RECT 6.96 3.8 7.44 7.92 ;
			RECT 6.96 5.42 7.6 7.92 ;
			RECT 1.24 7.44 7.6 7.92 ;
			RECT 1.24 7.44 1.72 8.94 ;
			RECT 1.08 8.3 1.72 8.94 ;
			RECT 6 7.44 6.64 10.08 ;
			RECT 4.6 8.44 5.24 11.1 ;
			RECT 7.44 10.46 8.08 11.1 ;
			RECT 4.6 10.62 8.08 11.1 ;
			RECT 9.24 2.18 9.88 3.5 ;
			RECT 8.12 3.02 9.88 3.5 ;
			RECT 8.12 3.02 8.6 9.94 ;
			RECT 8.12 9.46 11.2 9.94 ;
			RECT 10.56 9.46 11.2 10.1 ;
			RECT 10.4 2.14 12.6 2.78 ;
			RECT 10.4 2.14 10.88 7.74 ;
			RECT 9.12 7.26 10.88 7.74 ;
			RECT 9.12 7.26 9.76 8.94 ;

	END

END SCHMTTE

MACRO SCHMTT50E
	CLASS CORE ;
	FOREIGN SCHMTT50E 0 0  ;
	ORIGIN 0 0 ;
	SIZE 15.84 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.16 4.9 5.8 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 3.226 LAYER MTL1  ;
	END A
	PIN EN
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.88 6.28 2.52 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.267 LAYER MTL1  ;
	END EN
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 13.4 7.98 15.44 8.46 ;
			RECT 14.8 1.98 15.44 8.46 ;
			RECT 13.4 7.98 14.04 10.62 ;

		END 

		ANTENNADIFFAREA 4.467 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 15.84 13.68 ;
			RECT 14.8 8.98 15.44 13.68 ;
			RECT 12.4 4.3 13.12 5.94 ;
			RECT 12.4 4.3 12.88 10.02 ;
			RECT 12 9.54 12.64 13.68 ;
			RECT 2.88 8.44 3.52 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 15.84 1.46 ;
			RECT 11.4 3.3 14 3.78 ;
			RECT 13.36 -0.48 14 3.78 ;
			RECT 11.08 8.26 11.88 8.9 ;
			RECT 11.4 3.3 11.88 8.9 ;
			RECT 0.6 -0.48 1.24 4.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 6.04 3.74 6.96 4.38 ;
			RECT 6.48 3.74 6.96 5.9 ;
			RECT 6.96 5.42 7.6 7.92 ;
			RECT 1.4 7.44 7.6 7.92 ;
			RECT 1.4 7.44 1.88 8.94 ;
			RECT 1.24 8.3 1.88 8.94 ;
			RECT 6.16 7.44 6.8 10.08 ;
			RECT 4.8 2.74 8.12 3.22 ;
			RECT 4.8 2.74 5.28 4.38 ;
			RECT 4.64 3.74 5.28 4.38 ;
			RECT 7.48 2.74 8.12 4.46 ;
			RECT 4.76 8.44 5.4 11.1 ;
			RECT 7.6 10.46 8.24 11.1 ;
			RECT 4.76 10.62 8.24 11.1 ;
			RECT 9.24 2.82 9.88 5.5 ;
			RECT 8.12 5.02 9.88 5.5 ;
			RECT 8.12 5.02 8.6 9.94 ;
			RECT 8.12 9.46 11.2 9.94 ;
			RECT 10.56 9.46 11.2 10.1 ;
			RECT 10.4 2.14 12.6 2.78 ;
			RECT 10.4 2.14 10.88 7.74 ;
			RECT 9.12 7.26 10.88 7.74 ;
			RECT 9.12 7.26 9.76 8.94 ;

	END

END SCHMTT50E

MACRO SCHMTT50
	CLASS CORE ;
	FOREIGN SCHMTT50 0 0  ;
	ORIGIN 0 0 ;
	SIZE 12.96 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 3.96 1.04 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 3.629 LAYER MTL1  ;
	END A
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 11.92 1.98 12.56 11.22 ;
			RECT 10.4 1.98 12.56 4.06 ;

		END 

		ANTENNADIFFAREA 5.491 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 12.96 13.68 ;
			RECT 10.04 5.42 10.68 10.66 ;
			RECT 9.68 10.14 10.32 13.68 ;
			RECT 0.4 10.46 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 12.96 1.46 ;
			RECT 8.8 -0.48 9.6 3.98 ;
			RECT 8.8 -0.48 9.44 9.62 ;
			RECT 1 -0.48 1.64 2.54 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 5.92 2.96 6.56 5.7 ;
			RECT 3.52 5.06 6.56 5.7 ;
			RECT 3.52 5.06 4.16 10.22 ;
			RECT 7.56 2.96 8.2 6.7 ;
			RECT 6.28 6.22 8.2 6.7 ;
			RECT 6.28 6.22 6.92 10.22 ;
			RECT 2.52 3.34 3.72 3.98 ;
			RECT 2.52 3.34 3 11.22 ;
			RECT 8.28 10.14 8.92 11.22 ;
			RECT 2.52 10.74 8.92 11.22 ;

	END

END SCHMTT50

MACRO SCHMTT25E
	CLASS CORE ;
	FOREIGN SCHMTT25E 0 0  ;
	ORIGIN 0 0 ;
	SIZE 15.84 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.92 4.9 5.56 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 3.312 LAYER MTL1  ;
	END A
	PIN EN
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.88 6.28 2.52 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.267 LAYER MTL1  ;
	END EN
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 13.4 7.98 15.44 8.46 ;
			RECT 14.8 1.98 15.44 8.46 ;
			RECT 13.4 7.98 14.04 10.62 ;

		END 

		ANTENNADIFFAREA 4.467 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 15.84 13.68 ;
			RECT 14.8 8.98 15.44 13.68 ;
			RECT 12.4 4.3 13.12 5.94 ;
			RECT 12.4 4.3 12.88 10.02 ;
			RECT 12 9.54 12.64 13.68 ;
			RECT 2.88 8.44 3.52 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 15.84 1.46 ;
			RECT 11.4 3.3 14 3.78 ;
			RECT 13.36 -0.48 14 3.78 ;
			RECT 11.08 8.26 11.88 8.9 ;
			RECT 11.4 3.3 11.88 8.9 ;
			RECT 0.48 -0.48 1.12 4.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 5.8 3.74 6.6 4.38 ;
			RECT 6.12 3.74 6.6 5.9 ;
			RECT 6.12 5.42 7.6 5.9 ;
			RECT 6.96 5.42 7.6 7.92 ;
			RECT 1.4 7.44 7.6 7.92 ;
			RECT 1.4 7.44 1.88 8.94 ;
			RECT 1.24 8.3 1.88 8.94 ;
			RECT 6.16 7.44 6.8 10.08 ;
			RECT 4.56 2.74 7.88 3.22 ;
			RECT 4.56 2.74 5.04 4.38 ;
			RECT 4.4 3.74 5.04 4.38 ;
			RECT 7.24 2.74 7.88 4.54 ;
			RECT 4.76 8.44 5.4 11.1 ;
			RECT 7.6 10.46 8.24 11.1 ;
			RECT 4.76 10.62 8.24 11.1 ;
			RECT 9.24 3.9 9.88 5.54 ;
			RECT 8.12 5.06 9.88 5.54 ;
			RECT 8.12 5.06 8.6 9.94 ;
			RECT 8.12 9.46 11.2 9.94 ;
			RECT 10.56 9.46 11.2 10.1 ;
			RECT 10.4 2.14 12.6 2.78 ;
			RECT 10.4 2.14 10.88 7.74 ;
			RECT 9.12 7.26 10.88 7.74 ;
			RECT 9.12 7.26 9.76 8.94 ;

	END

END SCHMTT25E

MACRO SCHMTT25
	CLASS CORE ;
	FOREIGN SCHMTT25 0 0  ;
	ORIGIN 0 0 ;
	SIZE 12.96 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 3.96 1.04 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 3.629 LAYER MTL1  ;
	END A
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 11.36 8.22 12.56 11.22 ;
			RECT 11.92 1.98 12.56 11.22 ;
			RECT 10.76 1.98 12.56 4.06 ;

		END 

		ANTENNADIFFAREA 5.491 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 12.96 13.68 ;
			RECT 9.44 5.42 10.08 10.5 ;
			RECT 9.12 9.98 9.76 13.68 ;
			RECT 0.4 10.46 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 12.96 1.46 ;
			RECT 9.12 -0.48 9.96 4.06 ;
			RECT 8.44 4.26 9.6 4.78 ;
			RECT 9.12 -0.48 9.6 4.78 ;
			RECT 8.24 7.82 8.92 9.46 ;
			RECT 8.44 4.26 8.92 9.46 ;
			RECT 1 -0.48 1.64 2.54 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 6.28 1.98 6.92 5.7 ;
			RECT 3.52 5.06 6.92 5.7 ;
			RECT 3.52 5.06 4.16 10.22 ;
			RECT 2.52 3.34 3.6 3.98 ;
			RECT 2.52 3.34 3 11.22 ;
			RECT 7.72 10.14 8.36 11.22 ;
			RECT 2.52 10.74 8.36 11.22 ;
			RECT 7.44 2.96 8.56 3.6 ;
			RECT 7.44 2.96 7.92 6.7 ;
			RECT 6.28 6.22 7.92 6.7 ;
			RECT 6.28 6.22 6.92 10.22 ;

	END

END SCHMTT25

MACRO SCHMTT
	CLASS CORE ;
	FOREIGN SCHMTT 0 0  ;
	ORIGIN 0 0 ;
	SIZE 14.4 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 4.96 2.04 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 3.629 LAYER MTL1  ;
	END A
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 11.9 8.22 14 8.78 ;
			RECT 13.36 1.98 14 8.78 ;
			RECT 13.34 1.98 14 4.06 ;
			RECT 11.9 8.22 12.54 11.22 ;

		END 

		ANTENNADIFFAREA 5.352 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 14.4 13.68 ;
			RECT 13.24 9.58 14 13.68 ;
			RECT 10.2 6.22 11.84 6.86 ;
			RECT 10.5 10.54 11.16 13.68 ;
			RECT 10.68 6.22 11.16 13.68 ;
			RECT 0.58 8.96 1.22 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 14.4 1.46 ;
			RECT 11.86 -0.48 12.5 4.06 ;
			RECT 9.18 5.14 12.34 5.66 ;
			RECT 11.86 -0.48 12.34 5.66 ;
			RECT 9.18 7.98 9.82 9.62 ;
			RECT 9.18 5.14 9.66 9.62 ;
			RECT 4.82 -0.48 5.46 2.54 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 2.74 8.72 3.38 9.36 ;
			RECT 2.9 8.72 3.38 10.22 ;
			RECT 5.9 8.4 6.54 10.22 ;
			RECT 2.9 9.74 6.54 10.22 ;
			RECT 8.78 1.98 9.42 3.62 ;
			RECT 6.66 3.12 9.42 3.62 ;
			RECT 6.66 3.12 7.14 5.34 ;
			RECT 4.22 4.7 7.14 5.34 ;
			RECT 4.22 4.7 4.86 8.94 ;
			RECT 3.04 3.74 3.68 7.94 ;
			RECT 1.74 7.46 3.68 7.94 ;
			RECT 1.74 7.46 2.22 11.22 ;
			RECT 9.06 10.58 9.7 11.22 ;
			RECT 1.74 10.74 9.7 11.22 ;
			RECT 10.42 2.96 11.06 4.62 ;
			RECT 7.66 4.14 11.06 4.62 ;
			RECT 7.66 4.14 8.3 9.04 ;

	END

END SCHMTT

MACRO OR4XL
	CLASS CORE ;
	FOREIGN OR4XL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 8.64 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 6.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.123 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.96 2.48 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.123 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.28 3.92 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.123 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 7.6 5.36 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.123 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.34 10.58 8.24 11.22 ;
			RECT 7.6 2.54 8.24 11.22 ;

		END 

		ANTENNADIFFAREA 1.689 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 8.64 13.68 ;
			RECT 4.8 10.7 5.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 8.64 1.46 ;
			RECT 5.92 -0.48 6.56 3.18 ;
			RECT 2.56 -0.48 3.2 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 4.24 3.54 4.88 4.22 ;
			RECT 1 3.54 1.66 4.22 ;
			RECT 4.24 3.7 7.06 4.22 ;
			RECT 1 3.74 7.06 4.22 ;
			RECT 6.42 3.7 7.06 10.06 ;
			RECT 3.8 9.58 7.06 10.06 ;
			RECT 0.4 9.5 1.04 11.22 ;
			RECT 3.8 9.58 4.28 11.22 ;
			RECT 0.4 10.74 4.28 11.22 ;

	END

END OR4XL

MACRO OR4
	CLASS CORE ;
	FOREIGN OR4 0 0  ;
	ORIGIN 0 0 ;
	SIZE 8.64 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 3.64 1.04 4.28 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.555 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.96 2.48 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.555 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.22 3.92 7.86 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.555 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 4.96 5.36 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.555 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.98 9.44 8.24 11.22 ;
			RECT 7.6 1.98 8.24 11.22 ;

		END 

		ANTENNADIFFAREA 3.168 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 8.64 13.68 ;
			RECT 5.44 10.6 6.16 13.68 ;
			RECT 5.52 9.46 6.16 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 8.64 1.46 ;
			RECT 6.14 -0.48 6.78 2.62 ;
			RECT 3.28 -0.48 3.92 2.62 ;
			RECT 0.4 -0.48 1.04 2.62 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1.8 1.98 2.44 3.62 ;
			RECT 4.74 1.98 5.38 3.62 ;
			RECT 1.8 3.14 7.08 3.62 ;
			RECT 6.44 7.02 7.08 8.92 ;
			RECT 6.6 3.14 7.08 8.92 ;
			RECT 4.44 8.44 7.08 8.92 ;
			RECT 4.44 8.44 4.92 11.22 ;
			RECT 0.4 10.56 4.92 11.22 ;

	END

END OR4

MACRO OR3XL
	CLASS CORE ;
	FOREIGN OR3XL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 7.6 1.04 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.979 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 2.16 3.8 2.8 4.44 ;
			RECT 1.84 4.96 2.68 5.6 ;
			RECT 2.16 3.8 2.68 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.979 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.28 3.92 7.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.979 LAYER MTL1  ;
	END C
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 5.24 10.58 6.8 11.22 ;
			RECT 6.16 3.26 6.8 11.22 ;
			RECT 5.86 3.26 6.8 3.94 ;

		END 

		ANTENNADIFFAREA 1.614 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 3.8 10.34 4.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 4.86 -0.48 6.5 2.26 ;
			RECT 0.52 -0.48 2.16 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 3.22 1.98 3.86 3.26 ;
			RECT 1 2.78 5.34 3.26 ;
			RECT 1 2.78 1.64 3.9 ;
			RECT 4.7 2.78 5.34 4.64 ;
			RECT 4.8 2.78 5.34 9.82 ;
			RECT 4.8 9.18 5.44 9.82 ;
			RECT 0.4 9.34 5.44 9.82 ;
			RECT 0.4 9.34 1.04 11.22 ;

	END

END OR3XL

MACRO OR32AXL
	CLASS CORE ;
	FOREIGN OR32AXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 8.64 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 7.6 2.48 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.253 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 5.28 3.92 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.253 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 7.6 5.36 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.253 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 5.28 6.8 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.979 LAYER MTL1  ;
	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 7.6 8.24 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.979 LAYER MTL1  ;
	END E
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.58 8.76 8.24 11.22 ;
			RECT 0.4 8.76 8.24 9.24 ;
			RECT 0.4 4.16 4.04 4.64 ;
			RECT 3.4 3 4.04 4.64 ;
			RECT 0.4 8.76 2.38 11.22 ;
			RECT 0.4 3 1.24 3.64 ;
			RECT 0.4 3 1.04 11.22 ;
			RECT 0.38 7.6 1.04 8.24 ;

		END 

		ANTENNADIFFAREA 5.571 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 8.64 13.68 ;
			RECT 5.2 9.78 5.84 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 8.64 1.46 ;
			RECT 6.2 -0.48 6.84 3.64 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 2 1.98 5.44 2.46 ;
			RECT 2 1.98 2.64 3.64 ;
			RECT 4.8 1.98 5.44 4.68 ;
			RECT 7.6 2.98 8.24 4.68 ;
			RECT 4.8 4.16 8.24 4.68 ;

	END

END OR32AXL

MACRO OR32A
	CLASS CORE ;
	FOREIGN OR32A 0 0  ;
	ORIGIN 0 0 ;
	SIZE 14.4 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 3.64 2.48 4.28 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.779 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.24 4.96 4.88 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.779 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.6 6.28 8.24 6.94 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.779 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 9.04 4.96 9.68 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.261 LAYER MTL1  ;
	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 10.48 3.64 12.12 4.28 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.261 LAYER MTL1  ;
	END E
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 11.62 7.92 13.26 8.86 ;
			RECT 0.4 7.92 13.26 8.4 ;
			RECT 5.12 1.98 5.76 2.62 ;
			RECT 0.4 1.98 5.76 2.46 ;
			RECT 0.4 1.98 2.72 2.62 ;
			RECT 1.72 7.92 2.36 9.56 ;
			RECT 0.4 1.98 1.04 8.4 ;

		END 

		ANTENNADIFFAREA 9.406 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 14.4 13.68 ;
			RECT 9.54 10.62 11.18 13.68 ;
			RECT 6.88 10.32 7.52 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 14.4 1.46 ;
			RECT 7.92 -0.48 8.56 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 10.58 5.96 11.22 ;
			RECT 4.12 8.92 8.86 9.56 ;
			RECT 9.08 1.98 9.96 2.62 ;
			RECT 3.6 2.98 4.24 3.62 ;
			RECT 6.52 2.78 9.56 3.26 ;
			RECT 9.08 1.98 9.56 3.26 ;
			RECT 6.52 1.98 7.16 3.62 ;
			RECT 3.6 3.14 7.16 3.62 ;

	END

END OR32A

MACRO OR31AXL
	CLASS CORE ;
	FOREIGN OR31AXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.28 3.92 6.94 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.253 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.96 2.48 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.253 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 3.64 1.04 4.28 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.253 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 7.6 5.36 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.648 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.8 9.32 6.8 9.8 ;
			RECT 6.16 1.98 6.8 9.8 ;
			RECT 6.02 1.98 6.8 2.62 ;
			RECT 3.8 9.32 4.44 10.98 ;

		END 

		ANTENNADIFFAREA 3.365 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 5.32 10.5 5.96 13.68 ;
			RECT 0.4 8.66 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 3.22 -0.48 3.86 2.62 ;
			RECT 0.42 -0.48 1.06 2.62 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1.82 1.98 2.46 3.62 ;
			RECT 4.62 1.98 5.26 3.62 ;
			RECT 1.82 3.14 5.26 3.62 ;

	END

END OR31AXL

MACRO OR31A
	CLASS CORE ;
	FOREIGN OR31A 0 0  ;
	ORIGIN 0 0 ;
	SIZE 12.96 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.58 6.4 8.24 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.779 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 3.96 5.36 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.779 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 2.28 6.28 3.92 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.779 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 8.04 3.64 9.68 4.28 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.469 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 10.24 9.18 11.12 10.82 ;
			RECT 10.48 1.98 11.12 10.82 ;
			RECT 8.16 1.98 11.12 2.62 ;
			RECT 7.44 9.18 11.12 9.84 ;

		END 

		ANTENNADIFFAREA 7.224 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 12.96 13.68 ;
			RECT 11.68 9.54 12.32 13.68 ;
			RECT 1.8 9.7 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 12.96 1.46 ;
			RECT 5.36 -0.48 6 2.26 ;
			RECT 2.32 -0.48 2.96 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 8.7 6.64 9.18 ;
			RECT 3.2 8.7 6.64 9.4 ;
			RECT 6 8.7 6.64 10.06 ;
			RECT 0.4 8.7 1.04 11.22 ;
			RECT 3.2 8.7 3.86 11.22 ;
			RECT 3.84 1.98 4.48 3.26 ;
			RECT 6.76 1.98 7.4 3.26 ;
			RECT 3.84 2.78 7.4 3.26 ;
			RECT 4.6 9.92 5.24 11.22 ;
			RECT 4.6 10.58 9.48 11.22 ;

	END

END OR31A

MACRO OR3
	CLASS CORE ;
	FOREIGN OR3 0 0  ;
	ORIGIN 0 0 ;
	SIZE 8.64 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 6.28 1.04 7.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.325 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.96 3.2 5.6 ;
			RECT 2.48 3.96 3.2 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.325 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 3.96 5.36 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.325 LAYER MTL1  ;
	END C
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 5.24 9.44 8.24 11.22 ;
			RECT 7.6 1.98 8.24 11.22 ;
			RECT 6.88 1.98 8.24 2.66 ;

		END 

		ANTENNADIFFAREA 3.254 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 8.64 13.68 ;
			RECT 3.8 9.44 4.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 8.64 1.46 ;
			RECT 5.34 -0.48 5.98 2.26 ;
			RECT 2.06 -0.48 2.7 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.42 1.98 1.06 3.26 ;
			RECT 3.7 1.98 4.34 3.26 ;
			RECT 0.42 2.78 6.36 3.26 ;
			RECT 5.88 3.18 6.86 3.82 ;
			RECT 6.22 3.18 6.86 8.92 ;
			RECT 0.4 8.44 6.86 8.92 ;
			RECT 0.4 8.44 1.04 11.22 ;

	END

END OR3

MACRO OR2XL
	CLASS CORE ;
	FOREIGN OR2XL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 3.64 1.04 5.28 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.835 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 5.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.835 LAYER MTL1  ;
	END B
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 5.32 1.98 5.96 4.28 ;
			RECT 4.22 10.58 5.36 11.22 ;
			RECT 4.72 3.64 5.36 11.22 ;

		END 

		ANTENNADIFFAREA 1.845 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 2.82 10.58 3.46 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 3.68 -0.48 4.32 2.36 ;
			RECT 0.4 -0.48 1.04 2.36 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 2.04 1.98 2.68 3.36 ;
			RECT 2.04 2.88 4.2 3.36 ;
			RECT 3.56 2.88 4.2 10.06 ;
			RECT 0.4 9.58 4.2 10.06 ;
			RECT 0.4 9.58 1.04 10.9 ;

	END

END OR2XL

MACRO OR2N2AXL
	CLASS CORE ;
	FOREIGN OR2N2AXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 8.64 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 7.6 1.04 9.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.763 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.763 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 6.28 5.36 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.238 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 4.96 3.92 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.238 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 5.66 9.7 8.24 10.18 ;
			RECT 7.6 3.78 8.24 10.18 ;
			RECT 7.14 3.78 8.24 4.42 ;
			RECT 5.66 9.7 6.3 10.62 ;

		END 

		ANTENNADIFFAREA 3.472 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 8.64 13.68 ;
			RECT 7.14 10.7 7.78 13.68 ;
			RECT 3.22 10.7 3.86 13.68 ;
			RECT 0.4 10.7 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 8.64 1.46 ;
			RECT 5.72 -0.48 6.36 2.26 ;
			RECT 2.8 -0.48 3.44 2.62 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 1.98 2.28 2.62 ;
			RECT 1.8 1.98 2.28 3.62 ;
			RECT 1.8 3.14 4.2 3.62 ;
			RECT 3.72 3.14 4.2 4.36 ;
			RECT 3.72 3.88 6.58 4.36 ;
			RECT 6.1 4.94 6.9 6.58 ;
			RECT 6.1 3.88 6.58 9.18 ;
			RECT 4.54 8.7 6.58 9.18 ;
			RECT 4.54 8.7 5.02 10.18 ;
			RECT 1.8 9.7 5.02 10.18 ;
			RECT 1.8 9.7 2.44 11.22 ;
			RECT 4.2 1.98 5.2 2.62 ;
			RECT 4.72 1.98 5.2 3.26 ;
			RECT 7.16 1.98 7.8 3.26 ;
			RECT 4.72 2.78 7.8 3.26 ;

	END

END OR2N2AXL

MACRO OR2N2A
	CLASS CORE ;
	FOREIGN OR2N2A 0 0  ;
	ORIGIN 0 0 ;
	SIZE 10.08 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 7.6 1.04 9.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.763 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.763 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 6.28 6.8 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.462 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.72 4.96 5.36 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.462 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 9.44 9.68 10.02 ;
			RECT 9.04 1.98 9.68 10.02 ;
			RECT 8.46 1.98 9.68 2.64 ;
			RECT 7.6 9.44 8.28 11.08 ;

		END 

		ANTENNADIFFAREA 7.022 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 10.08 13.68 ;
			RECT 9.04 10.7 9.68 13.68 ;
			RECT 3.22 10.7 5.78 13.68 ;
			RECT 0.4 10.7 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 10.08 1.46 ;
			RECT 5.66 -0.48 6.3 2.36 ;
			RECT 2.82 -0.48 3.46 2.62 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 4.26 1.98 4.9 3.36 ;
			RECT 7.06 1.98 7.7 3.36 ;
			RECT 4.26 2.88 7.7 3.36 ;
			RECT 0.4 1.98 2.3 2.62 ;
			RECT 1.82 1.98 2.3 3.62 ;
			RECT 1.82 3.14 3.74 3.62 ;
			RECT 3.26 3.14 3.74 4.36 ;
			RECT 3.26 3.88 8.52 4.36 ;
			RECT 7.88 3.88 8.52 5.52 ;
			RECT 7.88 3.88 8.36 8.92 ;
			RECT 6.6 8.44 8.36 8.92 ;
			RECT 6.6 8.44 7.08 10.18 ;
			RECT 1.82 9.7 7.08 10.18 ;
			RECT 1.82 9.7 2.46 11.22 ;

	END

END OR2N2A

MACRO OR2N1AXL
	CLASS CORE ;
	FOREIGN OR2N1AXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 6.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.763 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 2.32 7.52 2.96 9.16 ;
			RECT 1.84 7.52 2.96 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.763 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 4.96 3.92 6.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.778 LAYER MTL1  ;
	END C
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.64 9.24 6.8 9.72 ;
			RECT 6.16 1.98 6.8 9.72 ;
			RECT 5.24 1.98 6.8 2.64 ;
			RECT 4.64 9.24 5.4 11.22 ;

		END 

		ANTENNADIFFAREA 2.131 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 6.04 10.7 6.68 13.68 ;
			RECT 3.2 10.68 3.84 13.68 ;
			RECT 0.4 10.7 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 2.82 -0.48 3.46 2.62 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 1.98 2.3 2.62 ;
			RECT 1.82 1.98 2.3 3.64 ;
			RECT 1.82 3.16 5.36 3.64 ;
			RECT 4.7 3.16 5.36 5.1 ;
			RECT 4.7 3.16 5.18 8.72 ;
			RECT 3.64 8.24 5.18 8.72 ;
			RECT 3.64 8.24 4.12 10.16 ;
			RECT 1.8 9.68 4.12 10.16 ;
			RECT 1.8 9.68 2.44 11.22 ;

	END

END OR2N1AXL

MACRO OR2N1A
	CLASS CORE ;
	FOREIGN OR2N1A 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 6.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.763 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 2.32 7.52 2.96 9.16 ;
			RECT 1.84 7.52 2.96 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.763 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 4.96 3.92 6.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.512 LAYER MTL1  ;
	END C
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.64 9.48 6.8 10.18 ;
			RECT 6.16 1.98 6.8 10.18 ;
			RECT 5.24 1.98 6.8 2.64 ;
			RECT 4.64 9.48 5.4 11.22 ;

		END 

		ANTENNADIFFAREA 4.138 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 6.04 10.7 6.68 13.68 ;
			RECT 3.2 10.68 3.84 13.68 ;
			RECT 0.4 10.7 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 2.82 -0.48 3.46 2.62 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 1.98 2.3 2.62 ;
			RECT 1.82 1.98 2.3 3.64 ;
			RECT 1.82 3.16 5.36 3.64 ;
			RECT 4.7 3.16 5.36 5.1 ;
			RECT 4.7 3.16 5.18 8.4 ;
			RECT 3.64 7.92 5.18 8.4 ;
			RECT 3.64 7.92 4.12 10.16 ;
			RECT 1.8 9.68 4.12 10.16 ;
			RECT 1.8 9.68 2.44 11.22 ;

	END

END OR2N1A

MACRO OR22AXL
	CLASS CORE ;
	FOREIGN OR22AXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 7.6 1.04 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.979 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.979 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 4.96 3.94 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.979 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 6.6 5.36 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.979 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 5.22 8.92 6.8 11.2 ;
			RECT 6.16 4.48 6.8 11.2 ;
			RECT 4.72 4.48 6.8 4.96 ;
			RECT 4.72 2.98 5.36 4.96 ;
			RECT 0.4 8.92 6.8 9.4 ;
			RECT 0.4 8.92 1.04 11.22 ;

		END 

		ANTENNADIFFAREA 4.309 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 2.82 9.92 3.46 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 1.8 -0.48 2.44 2.62 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 3.2 1.98 6.76 2.46 ;
			RECT 0.4 1.98 1.04 3.62 ;
			RECT 3.2 1.98 3.84 3.62 ;
			RECT 0.4 3.14 3.84 3.62 ;
			RECT 6.12 1.98 6.76 3.62 ;

	END

END OR22AXL

MACRO OR22A
	CLASS CORE ;
	FOREIGN OR22A 0 0  ;
	ORIGIN 0 0 ;
	SIZE 8.64 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.84 6.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.261 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 3.96 3.92 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.261 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 6.22 5.36 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.261 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 4.96 6.8 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.261 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 3.16 8.24 10.88 ;
			RECT 0.4 8.28 8.24 8.94 ;
			RECT 5.34 3.16 8.24 3.64 ;
			RECT 5.34 2.98 5.98 3.64 ;
			RECT 0.4 8.28 1.04 11.22 ;

		END 

		ANTENNADIFFAREA 10.494 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 8.64 13.68 ;
			RECT 2.82 10.7 5.86 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 8.64 1.46 ;
			RECT 2.24 -0.48 2.88 2.36 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 3.64 1.98 7.5 2.46 ;
			RECT 6.86 1.98 7.5 2.64 ;
			RECT 0.84 2.36 1.48 3.36 ;
			RECT 3.64 1.98 4.28 3.36 ;
			RECT 0.84 2.88 4.28 3.36 ;

	END

END OR22A

MACRO OR222AXL
	CLASS CORE ;
	FOREIGN OR222AXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 10.08 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.28 3.92 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.051 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.96 2.48 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.051 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 7.6 5.36 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.051 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 7.6 1.04 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.051 LAYER MTL1  ;
	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 4.96 8.24 5.62 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.051 LAYER MTL1  ;
	END E
	PIN F
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 6.28 6.8 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.051 LAYER MTL1  ;
	END F
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 8.26 8.9 9.68 11.06 ;
			RECT 9.04 3.94 9.68 11.06 ;
			RECT 7.56 3.94 9.68 4.42 ;
			RECT 4.86 8.9 9.68 9.38 ;
			RECT 7.56 2.98 8.2 4.42 ;
			RECT 3.42 10.02 5.34 10.66 ;
			RECT 4.86 8.9 5.34 10.66 ;

		END 

		ANTENNADIFFAREA 5.23 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 10.08 13.68 ;
			RECT 5.86 9.9 6.5 13.68 ;
			RECT 1 8.78 1.64 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 10.08 1.46 ;
			RECT 3.16 -0.48 3.84 2.44 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1.8 1.98 2.44 3.44 ;
			RECT 4.6 1.98 5.24 3.44 ;
			RECT 1.8 2.96 5.24 3.44 ;
			RECT 6.14 1.98 9.62 2.46 ;
			RECT 0.4 1.98 1.04 2.64 ;
			RECT 8.98 1.98 9.62 3.42 ;
			RECT 0.56 1.98 1.04 4.44 ;
			RECT 6.14 1.98 6.78 4.44 ;
			RECT 0.56 3.96 6.78 4.44 ;

	END

END OR222AXL

MACRO OR222A
	CLASS CORE ;
	FOREIGN OR222A 0 0  ;
	ORIGIN 0 0 ;
	SIZE 12.96 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.84 6.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.376 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 4.86 4.92 5.5 ;
			RECT 3.28 4.86 3.92 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.376 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 5.16 6.22 6.8 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.376 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 4.96 8.24 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.376 LAYER MTL1  ;
	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 9.04 6.28 9.68 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.376 LAYER MTL1  ;
	END E
	PIN F
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 10.48 4.96 11.12 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.376 LAYER MTL1  ;
	END F
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 9.7 12.56 10.18 ;
			RECT 11.92 3.16 12.56 10.18 ;
			RECT 6.22 9.54 12.56 10.18 ;
			RECT 9.62 3.16 12.56 3.64 ;
			RECT 9.62 2.98 10.26 3.64 ;
			RECT 6.22 8.3 8.86 10.18 ;
			RECT 0.4 8.28 1.04 11.22 ;

		END 

		ANTENNADIFFAREA 11.04 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 12.96 13.68 ;
			RECT 9.76 10.7 11.4 13.68 ;
			RECT 2.82 10.7 5.86 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 12.96 1.46 ;
			RECT 2.24 -0.48 2.88 2.36 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.84 1.98 1.48 3.64 ;
			RECT 3.64 1.98 4.28 3.64 ;
			RECT 6.82 2.98 7.46 3.64 ;
			RECT 0.84 3.16 7.46 3.64 ;
			RECT 5.42 1.98 11.66 2.46 ;
			RECT 11.02 1.98 11.66 2.62 ;
			RECT 5.42 1.98 6.06 2.64 ;
			RECT 8.22 1.98 8.86 3.64 ;

	END

END OR222A

MACRO OR221AXL
	CLASS CORE ;
	FOREIGN OR221AXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 10.08 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.051 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 7.6 3.92 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.051 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 4.96 6.8 6.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.051 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 5.22 5.36 6.86 ;
			RECT 0.4 4.96 5.2 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.051 LAYER MTL1  ;
	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 7.6 8.24 9.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.72 LAYER MTL1  ;
	END E
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.82 10.74 9.68 11.22 ;
			RECT 9.04 2.68 9.68 11.22 ;
			RECT 8.04 10.58 9.68 11.22 ;
			RECT 7.64 2.68 9.68 3.34 ;
			RECT 3.82 10.58 4.54 11.22 ;

		END 

		ANTENNADIFFAREA 4.04 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 10.08 13.68 ;
			RECT 6.22 9.5 6.86 10.14 ;
			RECT 1.32 9.58 6.86 10.06 ;
			RECT 1.32 9.48 1.96 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 10.08 1.46 ;
			RECT 3.32 -0.48 3.96 2.36 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1.8 2.72 2.44 3.36 ;
			RECT 4.84 2.7 5.48 3.36 ;
			RECT 1.8 2.88 5.48 3.36 ;
			RECT 0.4 2.68 1.04 4.36 ;
			RECT 6.24 2.68 6.88 4.36 ;
			RECT 0.4 3.88 6.88 4.36 ;

	END

END OR221AXL

MACRO OR221A
	CLASS CORE ;
	FOREIGN OR221A 0 0  ;
	ORIGIN 0 0 ;
	SIZE 10.08 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.376 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.22 3.92 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.376 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 4.96 6.8 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.376 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.68 4.88 5.32 6.86 ;
			RECT 0.4 4.88 5.32 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.376 LAYER MTL1  ;
	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 6.14 8.24 7.78 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.584 LAYER MTL1  ;
	END E
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 2.8 10.58 9.68 11.22 ;
			RECT 9.04 2.4 9.68 11.22 ;
			RECT 7.4 2.4 9.68 3.06 ;

		END 

		ANTENNADIFFAREA 8.323 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 10.08 13.68 ;
			RECT 6.22 8.3 7.86 8.94 ;
			RECT 0.4 9.58 6.7 10.06 ;
			RECT 6.22 8.3 6.7 10.06 ;
			RECT 0.4 8.44 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 10.08 1.46 ;
			RECT 3.2 -0.48 3.84 2.36 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1.8 2.4 2.44 3.36 ;
			RECT 4.6 2.38 5.24 3.36 ;
			RECT 1.8 2.88 5.24 3.36 ;
			RECT 0.4 2.4 1.04 4.36 ;
			RECT 6 2.4 6.64 4.36 ;
			RECT 0.4 3.88 6.64 4.36 ;

	END

END OR221A

MACRO OR21AXL
	CLASS CORE ;
	FOREIGN OR21AXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 5.76 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 7.6 1.04 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.979 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.96 2.48 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.979 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.28 3.92 7.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.648 LAYER MTL1  ;
	END C
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.24 9.4 5.36 11.22 ;
			RECT 4.72 1.98 5.36 11.22 ;
			RECT 4.6 1.98 5.36 2.64 ;
			RECT 0.4 9.4 5.36 9.88 ;
			RECT 0.4 9.4 1.04 11.22 ;

		END 

		ANTENNADIFFAREA 3.344 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 5.76 13.68 ;
			RECT 2.8 10.4 3.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 5.76 1.46 ;
			RECT 1.8 -0.48 2.44 2.62 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 1.98 1.04 3.62 ;
			RECT 3.2 1.98 3.84 3.62 ;
			RECT 0.4 3.14 3.84 3.62 ;

	END

END OR21AXL

MACRO OR21A
	CLASS CORE ;
	FOREIGN OR21A 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.261 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 3.96 3.92 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.261 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 6.22 5.36 7.86 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.469 LAYER MTL1  ;
	END C
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 5.54 9.48 6.8 11.22 ;
			RECT 6.16 1.98 6.8 11.22 ;
			RECT 5.66 1.98 6.8 2.64 ;
			RECT 0.4 9.7 6.8 10.18 ;
			RECT 0.4 8.76 1.04 11.22 ;

		END 

		ANTENNADIFFAREA 7.59 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 2.82 10.7 3.46 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 2.82 -0.48 3.46 2.36 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1.36 1.98 2 3.36 ;
			RECT 4.26 1.98 4.9 3.36 ;
			RECT 1.36 2.88 4.9 3.36 ;

	END

END OR21A

MACRO OR211AXL
	CLASS CORE ;
	FOREIGN OR211AXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 3.96 1.04 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.051 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.051 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 7.6 3.94 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.72 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 5.28 5.36 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.72 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 5.66 9.54 6.8 11.22 ;
			RECT 6.16 1.98 6.8 11.22 ;
			RECT 5.66 1.98 6.8 2.62 ;
			RECT 2.82 9.54 6.8 10.04 ;
			RECT 2.82 9.54 3.46 11.22 ;

		END 

		ANTENNADIFFAREA 3.662 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 4.26 10.56 4.9 13.68 ;
			RECT 0.4 9.34 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 1.8 -0.48 2.44 2.42 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 1.98 1.04 3.42 ;
			RECT 3.2 1.98 3.84 3.42 ;
			RECT 0.4 2.94 3.84 3.42 ;

	END

END OR211AXL

MACRO OR211A
	CLASS CORE ;
	FOREIGN OR211A 0 0  ;
	ORIGIN 0 0 ;
	SIZE 8.64 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.84 6.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.376 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 4.96 3.92 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.376 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 6.28 5.36 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.584 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 7.6 6.8 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.584 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.06 8.92 8.24 11.22 ;
			RECT 7.6 1.98 8.24 11.22 ;
			RECT 6.66 1.98 8.24 3.62 ;
			RECT 4.26 8.92 8.24 9.42 ;
			RECT 2.82 10.58 4.9 11.22 ;
			RECT 4.26 8.92 4.9 11.22 ;

		END 

		ANTENNADIFFAREA 8.744 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 8.64 13.68 ;
			RECT 5.66 9.94 6.3 13.68 ;
			RECT 0.4 8.58 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 8.64 1.46 ;
			RECT 2.82 -0.48 3.46 2.62 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1.36 1.98 2 3.62 ;
			RECT 4.26 1.98 4.9 3.62 ;
			RECT 1.36 3.14 4.9 3.62 ;

	END

END OR211A

MACRO OR2
	CLASS CORE ;
	FOREIGN OR2 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 3.64 1.04 5.28 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.123 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 5.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.123 LAYER MTL1  ;
	END B
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.88 1.98 5.72 2.62 ;
			RECT 4.46 9.58 5.36 11.22 ;
			RECT 4.88 1.98 5.36 11.22 ;
			RECT 4.72 3.64 5.36 11.22 ;

		END 

		ANTENNADIFFAREA 3.194 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 2.94 9.76 3.58 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 3.68 -0.48 4.32 2.36 ;
			RECT 0.4 -0.48 1.04 2.36 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 2.04 1.98 2.68 3.36 ;
			RECT 2.04 2.88 4.1 3.36 ;
			RECT 3.46 2.88 4.1 7.92 ;
			RECT 3.46 2.88 3.94 9.24 ;
			RECT 0.4 8.76 3.94 9.24 ;
			RECT 0.4 8.76 1.04 11.22 ;

	END

END OR2

MACRO NOR5
	CLASS CORE ;
	FOREIGN NOR5 0 0  ;
	ORIGIN 0 0 ;
	SIZE 12.96 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 7.6 1.04 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.123 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.123 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 4.96 3.92 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.123 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 6.28 5.36 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.123 LAYER MTL1  ;
	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 3.96 6.8 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.123 LAYER MTL1  ;
	END E
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 10.48 3.64 12.56 4.12 ;
			RECT 11.92 1.98 12.56 4.12 ;
			RECT 10.48 9.02 11.36 11.22 ;
			RECT 10.48 3.64 11.12 11.22 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 12.96 13.68 ;
			RECT 9.32 9.02 9.96 13.68 ;
			RECT 6.24 9.92 6.88 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 12.96 1.46 ;
			RECT 10.52 -0.48 11.16 2.26 ;
			RECT 8.88 -0.48 9.52 2.26 ;
			RECT 4.8 -0.48 5.44 2.26 ;
			RECT 1 -0.48 1.64 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 3.16 1.98 3.8 3.26 ;
			RECT 6.44 1.98 7.08 3.26 ;
			RECT 1 2.78 7.8 3.26 ;
			RECT 1 2.78 1.64 3.9 ;
			RECT 7.32 3.98 8.44 5.62 ;
			RECT 7.32 2.78 7.8 9.4 ;
			RECT 5.24 8.92 7.8 9.4 ;
			RECT 0.84 9.18 1.48 11.22 ;
			RECT 5.24 8.92 5.72 11.22 ;
			RECT 0.84 10.74 5.72 11.22 ;
			RECT 8.96 3.26 9.72 3.9 ;
			RECT 8.96 3.26 9.44 8.5 ;
			RECT 8.32 7.86 9.96 8.5 ;
			RECT 8.32 7.86 8.8 11.14 ;
			RECT 7.76 10.5 8.8 11.14 ;

	END

END NOR5

MACRO NOR4XL
	CLASS CORE ;
	FOREIGN NOR4XL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.74 6.28 5.38 7.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.267 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 5.28 3.92 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.267 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.267 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.36 4.96 1 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.267 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.8 8.76 6.8 9.56 ;
			RECT 6.16 3.26 6.8 9.56 ;
			RECT 1.12 3.8 6.8 4.28 ;
			RECT 5.56 3.26 6.8 4.28 ;
			RECT 4.8 8.76 5.44 11.22 ;
			RECT 1.12 3.26 1.76 4.28 ;

		END 

		ANTENNADIFFAREA 4.8 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 0.4 8.76 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 5.56 -0.48 6.2 2.26 ;
			RECT 3.4 -0.48 4.04 3.28 ;
			RECT 1.12 -0.48 1.76 2.26 ;

		END 

	END gndd!

END NOR4XL

MACRO NOR4ANXL
	CLASS CORE ;
	FOREIGN NOR4ANXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 8.64 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 6.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.734 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 4.96 5.36 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.512 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.28 3.92 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.512 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.96 2.48 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.512 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 2.78 8.24 11.22 ;
			RECT 7 2.78 8.24 3.9 ;
			RECT 3.4 2.78 8.24 3.26 ;
			RECT 3.4 1.98 4.04 3.26 ;

		END 

		ANTENNADIFFAREA 5.132 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 8.64 13.68 ;
			RECT 1.86 10.74 2.5 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 8.64 1.46 ;
			RECT 7 -0.48 7.64 2.26 ;
			RECT 5.04 -0.48 5.68 2.26 ;
			RECT 1.7 -0.48 2.34 2.42 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1.18 3.44 1.82 4.26 ;
			RECT 1.18 3.78 6.46 4.26 ;
			RECT 5.98 5.42 7.08 7.06 ;
			RECT 5.98 3.78 6.46 9.18 ;
			RECT 0.4 8.7 6.46 9.18 ;
			RECT 0.4 8.7 1.04 9.34 ;

	END

END NOR4ANXL

MACRO NOR4
	CLASS CORE ;
	FOREIGN NOR4 0 0  ;
	ORIGIN 0 0 ;
	SIZE 12.96 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 6.28 9.24 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.707 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 4.02 6.8 5.66 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.707 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 3.8 4.92 4.44 ;
			RECT 3.28 3.64 3.92 4.44 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.707 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.84 2.32 2.48 2.96 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.707 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 10.6 7.92 11.24 9.82 ;
			RECT 10.48 2.78 11.12 8.66 ;
			RECT 4.64 2.78 11.12 3.26 ;
			RECT 7.56 1.98 8.2 3.26 ;
			RECT 4.64 1.98 5.28 3.26 ;

		END 

		ANTENNADIFFAREA 5.04 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 12.96 13.68 ;
			RECT 1.72 9.18 2.36 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 12.96 1.46 ;
			RECT 8.96 -0.48 9.6 2.26 ;
			RECT 6.16 -0.48 6.8 2.26 ;
			RECT 3.12 -0.48 3.76 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 8.18 3.56 8.66 ;
			RECT 2.92 8.18 3.56 11.22 ;
			RECT 0.4 8.18 1.04 11.22 ;
			RECT 2.92 10.58 5.96 11.22 ;
			RECT 4.12 9.18 8.84 9.82 ;
			RECT 7 10.58 12.44 11.22 ;

	END

END NOR4

MACRO NOR3XL
	CLASS CORE ;
	FOREIGN NOR3XL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 5.76 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 7.6 3.92 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.181 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.181 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 4.96 1.04 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.181 LAYER MTL1  ;
	END C
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.8 8.92 5.36 10.88 ;
			RECT 4.72 3.64 5.36 10.88 ;
			RECT 1.4 3.96 5.36 4.44 ;
			RECT 4.68 3.64 5.36 4.44 ;
			RECT 1.4 3.78 2.04 4.44 ;

		END 

		ANTENNADIFFAREA 4.173 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 5.76 13.68 ;
			RECT 0.4 8.7 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 5.76 1.46 ;
			RECT 3.04 -0.48 3.68 3.44 ;
			RECT 1.4 -0.48 2.04 2.26 ;

		END 

	END gndd!

END NOR3XL

MACRO NOR3ANXL
	CLASS CORE ;
	FOREIGN NOR3ANXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 8.92 1.04 9.56 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.691 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 5.28 3.92 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.181 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 7.6 2.48 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.181 LAYER MTL1  ;
	END C
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 2.86 6.8 11.22 ;
			RECT 3.16 2.86 6.8 3.34 ;
			RECT 3.16 1.98 3.8 3.34 ;

		END 

		ANTENNADIFFAREA 4.363 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 2.72 10.7 3.36 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 5.6 -0.48 6.24 2.34 ;
			RECT 1 -0.48 1.64 2.34 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1 3.34 1.66 3.98 ;
			RECT 1.12 3.86 5.46 4.38 ;
			RECT 4.98 4.34 5.62 5.98 ;
			RECT 4.98 3.86 5.46 10.18 ;
			RECT 1.72 9.7 5.46 10.18 ;
			RECT 1.72 9.7 2.2 11.2 ;
			RECT 1.28 10.56 2.2 11.2 ;

	END

END NOR3ANXL

MACRO NOR3AN
	CLASS CORE ;
	FOREIGN NOR3AN 0 0  ;
	ORIGIN 0 0 ;
	SIZE 11.52 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 7.6 2.48 9.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.734 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 4.96 6.36 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.304 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.28 3.92 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.304 LAYER MTL1  ;
	END C
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.88 8.22 9.68 8.86 ;
			RECT 9.04 1.98 9.68 8.86 ;
			RECT 4.38 2.86 9.68 3.34 ;
			RECT 7.32 1.98 9.68 3.34 ;
			RECT 7.66 8.22 8.3 10.88 ;
			RECT 4.38 1.98 5.02 3.34 ;

		END 

		ANTENNADIFFAREA 6.929 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 11.52 13.68 ;
			RECT 2.9 10.76 3.54 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 11.52 1.46 ;
			RECT 5.92 -0.48 6.56 2.34 ;
			RECT 2.84 -0.48 3.48 2.34 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1.2 1.98 1.84 2.62 ;
			RECT 1.32 1.98 1.84 3.4 ;
			RECT 1.32 2.92 3.86 3.4 ;
			RECT 3.38 2.92 3.86 4.34 ;
			RECT 3.38 3.86 7.54 4.34 ;
			RECT 7.04 3.86 7.54 7.7 ;
			RECT 5.88 7.06 7.54 7.7 ;
			RECT 5.88 7.06 6.36 10.24 ;
			RECT 1.54 9.76 6.36 10.24 ;
			RECT 1.54 9.76 2.02 11.2 ;
			RECT 1.38 10.56 2.02 11.2 ;

	END

END NOR3AN

MACRO NOR3
	CLASS CORE ;
	FOREIGN NOR3 0 0  ;
	ORIGIN 0 0 ;
	SIZE 11.52 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.6 6.28 8.24 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.347 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 3.96 5.36 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.347 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 2.28 6.28 3.92 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.347 LAYER MTL1  ;
	END C
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 8.28 8.22 9.68 11.22 ;
			RECT 9.04 1.98 9.68 11.22 ;
			RECT 4.38 2.86 9.68 3.34 ;
			RECT 7.32 1.98 9.68 3.34 ;
			RECT 7.28 8.22 9.68 8.86 ;
			RECT 4.38 1.98 5.02 3.34 ;

		END 

		ANTENNADIFFAREA 7.297 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 11.52 13.68 ;
			RECT 3.52 8.7 4.16 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 11.52 1.46 ;
			RECT 5.92 -0.48 6.56 2.34 ;
			RECT 2.84 -0.48 3.48 2.34 ;

		END 

	END gndd!

END NOR3

MACRO NOR2XL
	CLASS CORE ;
	FOREIGN NOR2XL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 4.32 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.907 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 7.6 1.04 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.907 LAYER MTL1  ;
	END B
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 2.8 9.4 3.92 11.22 ;
			RECT 3.28 3.26 3.92 11.22 ;
			RECT 2.68 3.26 3.92 3.9 ;

		END 

		ANTENNADIFFAREA 2.84 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 4.32 13.68 ;
			RECT 0.4 9.7 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 4.32 1.46 ;
			RECT 2.92 -0.48 3.56 2.26 ;
			RECT 0.52 -0.48 1.16 2.9 ;

		END 

	END gndd!

END NOR2XL

MACRO NOR2ANXL
	CLASS CORE ;
	FOREIGN NOR2ANXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 5.76 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 7.54 1.04 9.18 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.734 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.96 2.48 6.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.138 LAYER MTL1  ;
	END B
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.24 8.92 5.36 11.22 ;
			RECT 4.72 2.32 5.36 11.22 ;
			RECT 4 3.1 5.36 3.74 ;

		END 

		ANTENNADIFFAREA 3.419 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 5.76 13.68 ;
			RECT 1.84 10.7 2.48 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 5.76 1.46 ;
			RECT 2.04 -0.48 2.68 2.3 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 2.78 1.04 3.42 ;
			RECT 0.4 2.94 3.48 3.42 ;
			RECT 3 5.78 4.04 7.42 ;
			RECT 3 2.94 3.48 10.18 ;
			RECT 0.84 9.7 3.48 10.18 ;
			RECT 0.84 9.7 1.32 11.1 ;
			RECT 0.4 10.42 1.32 11.1 ;

	END

END NOR2ANXL

MACRO NOR2AN
	CLASS CORE ;
	FOREIGN NOR2AN 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 6.28 1.04 7.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.734 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.02 2.48 5.66 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.304 LAYER MTL1  ;
	END B
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.28 8.4 6.8 9.56 ;
			RECT 4.88 2 5.36 9.56 ;
			RECT 4.72 2 5.36 5.6 ;

		END 

		ANTENNADIFFAREA 6.007 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 1.84 10.9 4.44 13.68 ;
			RECT 1.84 9.9 2.48 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 6.12 -0.48 6.76 2.36 ;
			RECT 3.32 -0.48 3.96 2.36 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1.66 1.98 2.3 3.36 ;
			RECT 1.66 2.88 4.2 3.36 ;
			RECT 3.72 2.88 4.2 7.86 ;
			RECT 3.72 6.22 4.36 7.86 ;
			RECT 3.28 7.34 3.76 9.24 ;
			RECT 0.84 8.76 3.76 9.24 ;
			RECT 0.84 8.76 1.32 11.1 ;
			RECT 0.4 10.42 1.32 11.1 ;

	END

END NOR2AN

MACRO NOR2
	CLASS CORE ;
	FOREIGN NOR2 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 4.96 3.92 6.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.059 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 2.64 2.48 4.28 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.059 LAYER MTL1  ;
	END B
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.56 9.58 5.36 10.22 ;
			RECT 4.72 2.12 5.36 10.22 ;

		END 

		ANTENNADIFFAREA 3.557 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 1.8 9.8 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 6.12 -0.48 6.76 2.36 ;
			RECT 3.32 -0.48 3.96 2.36 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 8.76 3.84 9.28 ;
			RECT 3.2 8.76 3.84 11.22 ;
			RECT 0.4 8.76 1.04 11.22 ;
			RECT 6 9.12 6.64 11.22 ;
			RECT 3.2 10.74 6.64 11.22 ;

	END

END NOR2

MACRO NAND7
	CLASS CORE ;
	FOREIGN NAND7 0 0  ;
	ORIGIN 0 0 ;
	SIZE 15.84 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 8.92 1.04 9.56 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.864 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.96 2.48 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.864 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 7.6 3.92 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.864 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 6.28 5.36 7.06 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.864 LAYER MTL1  ;
	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 7.6 6.8 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.864 LAYER MTL1  ;
	END E
	PIN F
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 6.28 8.24 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.864 LAYER MTL1  ;
	END F
	PIN G
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 9.04 4.96 9.68 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.864 LAYER MTL1  ;
	END G
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 14.56 8.02 15.2 11.22 ;
			RECT 13.36 8.02 15.2 8.5 ;
			RECT 13.36 1.98 14 8.5 ;
			RECT 12.72 1.98 14 2.62 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 15.84 13.68 ;
			RECT 13.16 9.02 13.8 13.68 ;
			RECT 8.8 10.7 9.44 13.68 ;
			RECT 6 10.7 6.64 13.68 ;
			RECT 3.2 10.7 3.84 13.68 ;
			RECT 0.4 10.7 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 15.84 1.46 ;
			RECT 11.32 -0.48 11.96 2.26 ;
			RECT 7.8 -0.48 8.44 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 1.98 7.28 2.62 ;
			RECT 6.8 1.98 7.28 3.26 ;
			RECT 6.8 2.78 8.92 3.26 ;
			RECT 8.44 2.78 8.92 4.26 ;
			RECT 8.44 3.78 11.08 4.26 ;
			RECT 1.8 9.7 11.08 10.18 ;
			RECT 1.8 9.7 2.44 11.22 ;
			RECT 4.6 9.7 5.24 11.22 ;
			RECT 7.4 9.7 8.04 11.22 ;
			RECT 10.44 3.78 11.08 11.22 ;
			RECT 10.2 9.7 11.08 11.22 ;
			RECT 9.44 1.98 10.08 3.26 ;
			RECT 9.44 2.78 12.2 3.26 ;
			RECT 11.64 3.14 12.84 4.78 ;
			RECT 11.64 3.14 12.28 10.88 ;

	END

END NAND7

MACRO NAND6
	CLASS CORE ;
	FOREIGN NAND6 0 0  ;
	ORIGIN 0 0 ;
	SIZE 14.4 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 8.92 1.04 9.56 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.864 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.96 2.48 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.864 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 7.6 3.92 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.864 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 6.28 5.36 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.864 LAYER MTL1  ;
	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 7.6 6.8 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.864 LAYER MTL1  ;
	END E
	PIN F
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 6.28 8.24 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.864 LAYER MTL1  ;
	END F
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 11.92 1.98 12.56 11.22 ;
			RECT 11.28 1.98 12.56 2.62 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 14.4 13.68 ;
			RECT 13.32 9.02 13.96 13.68 ;
			RECT 8.8 10.7 9.44 13.68 ;
			RECT 6 10.7 6.64 13.68 ;
			RECT 3.2 10.7 3.84 13.68 ;
			RECT 0.4 10.7 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 14.4 1.46 ;
			RECT 9.88 -0.48 10.52 2.26 ;
			RECT 6.8 -0.48 7.44 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 1.98 6.28 2.62 ;
			RECT 5.8 1.98 6.28 3.26 ;
			RECT 5.8 2.78 7.92 3.26 ;
			RECT 7.44 2.78 7.92 4.26 ;
			RECT 7.44 3.78 9.4 4.26 ;
			RECT 8.76 3.78 9.4 10.18 ;
			RECT 1.8 9.7 9.4 10.18 ;
			RECT 1.8 9.7 2.44 11.22 ;
			RECT 4.6 9.7 5.24 11.22 ;
			RECT 7.4 9.7 8.04 11.22 ;
			RECT 8.44 1.98 9.08 3.26 ;
			RECT 8.44 2.78 10.44 3.26 ;
			RECT 9.92 3.14 11.4 4.78 ;
			RECT 9.92 2.78 10.4 10.18 ;
			RECT 10.32 9.7 10.96 10.86 ;

	END

END NAND6

MACRO NAND5
	CLASS CORE ;
	FOREIGN NAND5 0 0  ;
	ORIGIN 0 0 ;
	SIZE 8.64 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.96 2.48 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.958 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3 6.28 3.92 6.92 ;
			RECT 2.92 7.28 3.56 7.92 ;
			RECT 3 6.28 3.56 7.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.958 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 6.28 5.36 7.62 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.958 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 6.28 6.8 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.958 LAYER MTL1  ;
	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 4.96 8.24 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.958 LAYER MTL1  ;
	END E
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 8.62 8.24 11.22 ;
			RECT 0.4 8.62 8.24 9.1 ;
			RECT 4.8 8.62 5.44 11.22 ;
			RECT 2 8.62 2.64 11.22 ;
			RECT 0.4 1.98 2.4 4.44 ;
			RECT 0.4 1.98 1.04 9.1 ;

		END 

		ANTENNADIFFAREA 9.862 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 8.64 13.68 ;
			RECT 6.2 9.62 6.84 13.68 ;
			RECT 3.4 9.62 4.04 13.68 ;
			RECT 0.6 9.62 1.24 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 8.64 1.46 ;
			RECT 7.16 -0.48 7.8 3.44 ;

		END 

	END gndd!

END NAND5

MACRO NAND4XL
	CLASS CORE ;
	FOREIGN NAND4XL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.96 2.48 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.749 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.28 3.92 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.749 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 7.6 5.36 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.749 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 8.92 6.8 9.56 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.749 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.76 9.7 5.4 11.22 ;
			RECT 0.4 9.7 5.4 10.18 ;
			RECT 1.96 9.7 2.6 11.22 ;
			RECT 0.4 1.98 2.4 2.62 ;
			RECT 0.4 1.98 1.04 10.18 ;

		END 

		ANTENNADIFFAREA 3.078 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 6.16 10.7 6.8 13.68 ;
			RECT 3.36 10.7 4 13.68 ;
			RECT 0.56 10.7 1.2 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 6.16 -0.48 6.8 2.62 ;

		END 

	END gndd!

END NAND4XL

MACRO NAND4ANXL
	CLASS CORE ;
	FOREIGN NAND4ANXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 8.64 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 3.64 8.24 4.28 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.691 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.28 3.92 8.06 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.85 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 6.28 5.36 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.85 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 4.96 6.8 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.85 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 9.7 5.36 11.22 ;
			RECT 0.4 9.7 5.36 10.18 ;
			RECT 1.8 9.7 2.44 11.22 ;
			RECT 0.4 1.98 1.66 2.62 ;
			RECT 0.4 1.98 1.04 10.18 ;

		END 

		ANTENNADIFFAREA 3.893 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 8.64 13.68 ;
			RECT 6.2 10.62 6.84 13.68 ;
			RECT 3.32 10.7 3.96 13.68 ;
			RECT 0.4 10.7 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 8.64 1.46 ;
			RECT 5.44 -0.48 6.08 2.3 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 6.6 1.98 7.72 2.62 ;
			RECT 2.18 2.84 7.08 3.32 ;
			RECT 6.6 1.98 7.08 3.32 ;
			RECT 1.56 3.14 2.66 3.62 ;
			RECT 1.56 3.14 2.2 5.04 ;
			RECT 1.56 3.14 2.04 9.18 ;
			RECT 1.56 8.7 6.7 9.18 ;
			RECT 6.16 8.7 6.7 10.1 ;
			RECT 6.16 9.62 8.08 10.1 ;
			RECT 7.6 9.62 8.08 10.86 ;
			RECT 7.6 10.22 8.24 10.86 ;

	END

END NAND4ANXL

MACRO NAND4AN
	CLASS CORE ;
	FOREIGN NAND4AN 0 0  ;
	ORIGIN 0 0 ;
	SIZE 8.64 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 7.6 8.24 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.691 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.28 3.92 7.06 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.973 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 6.28 5.36 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.973 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 4.96 6.8 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.973 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 9.44 5.36 11.22 ;
			RECT 0.4 9.44 5.36 9.92 ;
			RECT 1.8 9.44 2.44 11.22 ;
			RECT 0.4 1.98 2.18 2.62 ;
			RECT 0.4 1.98 1.04 9.92 ;

		END 

		ANTENNADIFFAREA 8.902 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 8.64 13.68 ;
			RECT 6.2 10.02 6.84 13.68 ;
			RECT 3.32 10.44 3.96 13.68 ;
			RECT 0.4 10.44 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 8.64 1.46 ;
			RECT 5.96 -0.48 6.6 2.44 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 7.12 1.98 8.24 2.62 ;
			RECT 2.7 2.96 7.6 3.44 ;
			RECT 7.12 1.98 7.6 3.44 ;
			RECT 1.56 3.14 3.18 3.62 ;
			RECT 1.56 3.14 2.2 6.04 ;
			RECT 1.56 3.14 2.04 8.92 ;
			RECT 1.56 8.44 6.7 8.92 ;
			RECT 6.16 8.76 8.24 9.24 ;
			RECT 7.6 8.76 8.24 10.86 ;

	END

END NAND4AN

MACRO NAND42
	CLASS CORE ;
	FOREIGN NAND42 0 0  ;
	ORIGIN 0 0 ;
	SIZE 14.4 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 5.3 2.48 6.94 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 3.542 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 5.28 5.36 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 3.542 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 5.28 8.24 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 3.542 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 10.48 6.28 12.12 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 3.542 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 10.2 8.7 10.84 11.22 ;
			RECT 0.4 8.7 10.84 9.18 ;
			RECT 7.4 8.7 8.04 11.22 ;
			RECT 4.6 8.7 5.24 11.22 ;
			RECT 1.8 8.7 2.44 11.22 ;
			RECT 0.4 4.28 2.44 4.76 ;
			RECT 1.8 2.98 2.44 4.76 ;
			RECT 0.4 4.28 1.04 9.18 ;

		END 

		ANTENNADIFFAREA 12.73 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 14.4 13.68 ;
			RECT 11.6 9.7 12.24 13.68 ;
			RECT 8.8 9.7 9.44 13.68 ;
			RECT 6 9.7 6.64 13.68 ;
			RECT 3.2 9.7 3.84 13.68 ;
			RECT 0.4 9.7 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 14.4 1.46 ;
			RECT 11.62 -0.48 12.32 3.76 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 1.98 6.64 2.46 ;
			RECT 0.4 1.98 1.04 3.76 ;
			RECT 6 1.98 6.64 3.76 ;
			RECT 3.2 1.98 3.84 4.02 ;
			RECT 4.6 2.98 5.24 4.76 ;
			RECT 8.84 2.98 9.48 4.76 ;
			RECT 4.6 4.28 9.48 4.76 ;
			RECT 7.44 1.98 10.88 2.46 ;
			RECT 7.44 1.98 8.08 3.76 ;
			RECT 10.24 1.98 10.88 4.76 ;
			RECT 13.04 1.98 13.68 4.76 ;
			RECT 10.24 4.28 13.68 4.76 ;

	END

END NAND42

MACRO NAND4
	CLASS CORE ;
	FOREIGN NAND4 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 5.14 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.771 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 5.98 3.92 7.62 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.771 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 6.28 5.36 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.771 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 4.96 6.8 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.771 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.76 8.62 5.4 11.22 ;
			RECT 0.4 8.62 5.4 9.1 ;
			RECT 1.96 8.62 2.6 11.22 ;
			RECT 0.4 1.98 2.4 3.64 ;
			RECT 0.4 1.98 1.04 9.1 ;

		END 

		ANTENNADIFFAREA 7.258 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 6.16 9.62 6.8 13.68 ;
			RECT 3.36 9.62 4 13.68 ;
			RECT 0.56 9.62 1.2 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 6.16 -0.48 6.8 3.26 ;

		END 

	END gndd!

END NAND4

MACRO NAND3XL
	CLASS CORE ;
	FOREIGN NAND3XL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 5.76 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 7.6 2.48 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.706 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.28 3.92 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.706 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 3.96 5.36 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.706 LAYER MTL1  ;
	END C
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 9.68 5.36 11.22 ;
			RECT 0.4 9.68 5.36 10.16 ;
			RECT 1.92 9.68 2.56 11.22 ;
			RECT 0.4 1.98 1.96 2.64 ;
			RECT 0.4 1.98 1.04 10.16 ;

		END 

		ANTENNADIFFAREA 2.806 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 5.76 13.68 ;
			RECT 3.32 10.68 3.96 13.68 ;
			RECT 0.52 10.68 1.16 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 5.76 1.46 ;
			RECT 4.72 -0.48 5.36 2.44 ;

		END 

	END gndd!

END NAND3XL

MACRO NAND3ANXL
	CLASS CORE ;
	FOREIGN NAND3ANXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 7.54 6.8 9.18 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.691 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 2.78 6.92 3.92 7.92 ;
			RECT 3.28 6.28 3.92 7.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.835 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.7 4.08 5.36 5.72 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.835 LAYER MTL1  ;
	END C
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.3 9.7 3.94 11.22 ;
			RECT 0.5 9.7 3.94 10.18 ;
			RECT 0.4 1.98 1.76 2.62 ;
			RECT 0.5 8.92 1.18 10.18 ;
			RECT 0.5 8.92 1.14 11.22 ;
			RECT 0.4 1.98 1.04 9.56 ;

		END 

		ANTENNADIFFAREA 3.498 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 4.74 10.7 5.38 13.68 ;
			RECT 1.9 10.7 2.54 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 4.52 -0.48 5.16 2.42 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 6.14 2.04 6.8 2.68 ;
			RECT 2.28 2.94 6.62 3.42 ;
			RECT 6.14 2.04 6.62 3.42 ;
			RECT 1.56 3.14 2.76 3.62 ;
			RECT 1.56 3.14 2.2 4.78 ;
			RECT 1.72 3.14 2.2 9.18 ;
			RECT 1.72 8.7 5.22 9.18 ;
			RECT 4.74 8.7 5.22 10.18 ;
			RECT 4.74 9.7 6.8 10.18 ;
			RECT 6.16 9.7 6.8 10.66 ;

	END

END NAND3ANXL

MACRO NAND3AN
	CLASS CORE ;
	FOREIGN NAND3AN 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 7.6 6.8 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.691 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.28 3.92 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.8 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 4.96 5.36 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.8 LAYER MTL1  ;
	END C
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.3 9.44 3.94 11.22 ;
			RECT 0.5 9.44 3.94 9.92 ;
			RECT 0.4 1.98 1.76 2.64 ;
			RECT 0.4 8.92 1.18 9.56 ;
			RECT 0.5 8.92 1.14 11.22 ;
			RECT 0.4 1.98 1.04 9.56 ;

		END 

		ANTENNADIFFAREA 7.52 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 4.74 10.02 5.38 13.68 ;
			RECT 1.9 10.44 2.54 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 4.52 -0.48 5.16 2.44 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 6.14 1.98 6.8 2.62 ;
			RECT 2.28 2.96 6.62 3.44 ;
			RECT 6.14 1.98 6.62 3.44 ;
			RECT 1.72 3.16 2.76 3.64 ;
			RECT 1.56 4 2.2 5.64 ;
			RECT 1.72 3.16 2.2 8.92 ;
			RECT 1.72 8.44 5.22 8.92 ;
			RECT 4.74 8.76 6.78 9.24 ;
			RECT 6.14 8.76 6.78 10.66 ;

	END

END NAND3AN

MACRO NAND32
	CLASS CORE ;
	FOREIGN NAND32 0 0  ;
	ORIGIN 0 0 ;
	SIZE 10.08 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.6 2.48 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 3.197 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.28 3.92 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 3.197 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 4.96 6.36 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 3.197 LAYER MTL1  ;
	END C
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.4 8.76 8.04 11.22 ;
			RECT 0.4 8.76 8.04 9.24 ;
			RECT 4.6 8.76 5.24 11.22 ;
			RECT 1.8 8.76 2.44 11.22 ;
			RECT 0.4 1.98 1.04 9.24 ;

		END 

		ANTENNADIFFAREA 11.053 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 10.08 13.68 ;
			RECT 8.8 9.22 9.44 13.68 ;
			RECT 5.98 10.08 6.64 13.68 ;
			RECT 3.2 10.08 3.84 13.68 ;
			RECT 0.4 10.08 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 10.08 1.46 ;
			RECT 5.8 -0.48 6.44 4.44 ;
			RECT 4.8 -0.48 6.44 2.26 ;

		END 

	END gndd!

END NAND32

MACRO NAND3
	CLASS CORE ;
	FOREIGN NAND3 0 0  ;
	ORIGIN 0 0 ;
	SIZE 5.76 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.96 2.48 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.598 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.28 3.92 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.598 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 7.6 5.36 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.598 LAYER MTL1  ;
	END C
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 8.94 5.36 11.22 ;
			RECT 0.4 8.94 5.36 9.42 ;
			RECT 1.92 8.94 2.56 11.22 ;
			RECT 0.4 1.98 1.96 3.64 ;
			RECT 0.4 1.98 1.04 9.56 ;

		END 

		ANTENNADIFFAREA 6.445 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 5.76 13.68 ;
			RECT 3.32 9.94 3.96 13.68 ;
			RECT 0.52 10.08 1.16 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 5.76 1.46 ;
			RECT 4.72 -0.48 5.36 3.36 ;

		END 

	END gndd!

END NAND3

MACRO NAND2XL
	CLASS CORE ;
	FOREIGN NAND2XL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 4.32 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 5.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.634 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 7.6 3.92 9.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.634 LAYER MTL1  ;
	END B
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.56 10.58 2.44 11.22 ;
			RECT 1.56 9.42 2.04 11.22 ;
			RECT 0.4 9.42 2.04 9.9 ;
			RECT 0.4 1.98 1.52 2.62 ;
			RECT 0.4 1.98 1.04 9.9 ;

		END 

		ANTENNADIFFAREA 1.715 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 4.32 13.68 ;
			RECT 3.2 10.66 3.84 13.68 ;
			RECT 0.4 10.66 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 4.32 1.46 ;
			RECT 3.28 -0.48 3.92 2.62 ;

		END 

	END gndd!

END NAND2XL

MACRO NAND2ANXL
	CLASS CORE ;
	FOREIGN NAND2ANXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 5.76 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 6.28 5.36 7.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.691 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 4 3.92 5.64 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.778 LAYER MTL1  ;
	END B
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.82 9.56 2.46 11.06 ;
			RECT 0.4 9.56 2.46 10.18 ;
			RECT 0.4 1.98 1.2 2.64 ;
			RECT 0.4 1.98 1.04 10.18 ;

		END 

		ANTENNADIFFAREA 2.218 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 5.76 13.68 ;
			RECT 3.32 10.7 3.96 13.68 ;
			RECT 0.42 10.7 1.06 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 5.76 1.46 ;
			RECT 3.08 -0.48 3.72 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 4.72 2 5.36 2.64 ;
			RECT 4.72 2 5.24 3.26 ;
			RECT 1.74 2.78 5.24 3.26 ;
			RECT 1.56 4 2.22 5.64 ;
			RECT 1.74 2.78 2.22 8.92 ;
			RECT 1.74 8.44 3.46 8.92 ;
			RECT 2.98 8.44 3.46 10.18 ;
			RECT 2.98 9.7 5.36 10.18 ;
			RECT 4.72 9.7 5.36 11.22 ;

	END

END NAND2ANXL

MACRO NAND2AN
	CLASS CORE ;
	FOREIGN NAND2AN 0 0  ;
	ORIGIN 0 0 ;
	SIZE 5.76 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 6.28 5.36 7.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.691 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 3.98 3.92 5.62 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.757 LAYER MTL1  ;
	END B
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.82 9.56 2.46 11.22 ;
			RECT 0.4 9.56 2.46 10.18 ;
			RECT 0.4 1.98 1.32 2.62 ;
			RECT 0.4 1.98 1.04 10.18 ;

		END 

		ANTENNADIFFAREA 4.998 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 5.76 13.68 ;
			RECT 3.32 10.64 3.96 13.68 ;
			RECT 0.42 10.7 1.06 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 5.76 1.46 ;
			RECT 3.08 -0.48 3.72 2.44 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 4.72 1.98 5.36 2.62 ;
			RECT 4.72 1.98 5.24 3.44 ;
			RECT 1.84 2.96 5.24 3.44 ;
			RECT 1.56 4.6 2.32 6.24 ;
			RECT 1.84 2.96 2.32 8.92 ;
			RECT 1.84 8.44 3.46 8.92 ;
			RECT 2.98 8.44 3.46 10.12 ;
			RECT 2.98 9.64 5.36 10.12 ;
			RECT 4.72 9.64 5.36 11.22 ;

	END

END NAND2AN

MACRO NAND22
	CLASS CORE ;
	FOREIGN NAND22 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 2.48 7.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.995 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.28 4.92 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.995 LAYER MTL1  ;
	END B
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.76 8.44 5.4 11.22 ;
			RECT 0.4 8.44 5.4 8.92 ;
			RECT 1.96 8.44 2.6 11.22 ;
			RECT 0.4 1.98 1.04 8.92 ;

		END 

		ANTENNADIFFAREA 8.086 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 6.16 9.5 6.8 13.68 ;
			RECT 3.36 9.44 4 13.68 ;
			RECT 0.56 9.5 1.2 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 3.16 -0.48 3.8 4.54 ;

		END 

	END gndd!

END NAND22

MACRO NAND2
	CLASS CORE ;
	FOREIGN NAND2 0 0  ;
	ORIGIN 0 0 ;
	SIZE 4.32 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.96 2.48 6.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.498 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.6 3.92 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.498 LAYER MTL1  ;
	END B
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.88 8.94 2.52 11.22 ;
			RECT 0.4 8.94 2.52 9.56 ;
			RECT 0.4 2.18 1.52 2.82 ;
			RECT 0.4 2.18 1.04 9.56 ;

		END 

		ANTENNADIFFAREA 4.058 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 4.32 13.68 ;
			RECT 3.28 9.7 3.92 13.68 ;
			RECT 0.48 10.08 1.12 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 4.32 1.46 ;
			RECT 3.28 -0.48 3.92 2.82 ;

		END 

	END gndd!

END NAND2

MACRO MUX41XL
	CLASS CORE ;
	FOREIGN MUX41XL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 25.92 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.562 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 4.14 6.8 9.34 ;
			RECT 6.04 4.14 6.8 4.78 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.562 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 4.14 8.24 9.34 ;
			RECT 7.4 4.14 8.24 4.78 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.562 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 12 2.84 12.64 3.48 ;
			RECT 11.92 3.64 12.56 9.34 ;
			RECT 12 2.84 12.56 9.34 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.562 LAYER MTL1  ;
	END D
	PIN S1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 13.32 8.7 14 9.34 ;
			RECT 13.36 4.2 14 9.34 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.685 LAYER MTL1  ;
	END S1
	PIN S2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 16.16 9.56 16.88 11.22 ;
			RECT 16.24 4.42 16.88 11.22 ;
			RECT 15.52 4.42 16.88 4.9 ;
			RECT 15.52 1.98 16 4.9 ;
			RECT 15.36 1.98 16 2.62 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.979 LAYER MTL1  ;
	END S2
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 24.88 3.64 25.52 11.02 ;
			RECT 24.28 3.64 25.52 4.28 ;

		END 

		ANTENNADIFFAREA 1.614 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 25.92 13.68 ;
			RECT 23.44 10.5 24.08 13.68 ;
			RECT 17.5 10.74 18.14 13.68 ;
			RECT 12.8 9.92 13.44 13.68 ;
			RECT 6.84 10.02 7.48 13.68 ;
			RECT 1.04 9.78 1.68 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 25.92 1.46 ;
			RECT 24.28 -0.48 24.92 2.64 ;
			RECT 16.52 -0.48 17.16 2.26 ;
			RECT 12.48 -0.48 13.12 2.28 ;
			RECT 6.4 -0.48 7.04 3.18 ;
			RECT 1 -0.48 1.64 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1.4 3.26 2.84 3.9 ;
			RECT 2.36 3.26 2.84 10.42 ;
			RECT 2.36 9.78 3.12 10.42 ;
			RECT 3.36 2.54 4.12 6.9 ;
			RECT 3.64 2.54 4.12 10.34 ;
			RECT 3.64 9.7 4.52 10.34 ;
			RECT 4.76 2.54 5.52 3.18 ;
			RECT 5.04 2.54 5.52 10.66 ;
			RECT 5.04 10.02 6.08 10.66 ;
			RECT 8.04 1.98 8.68 3.62 ;
			RECT 8.04 3.14 9.24 3.62 ;
			RECT 8.76 3.14 9.24 10.66 ;
			RECT 8.24 10.02 9.24 10.66 ;
			RECT 9.44 1.98 10.24 2.62 ;
			RECT 9.76 1.98 10.24 10.46 ;
			RECT 9.76 5.2 10.4 10.46 ;
			RECT 10.84 1.98 11.48 2.62 ;
			RECT 10.92 1.98 11.4 10.66 ;
			RECT 10.92 10.02 12.04 10.66 ;
			RECT 14.12 2.02 14.76 3.62 ;
			RECT 14.52 7.56 15.32 9.2 ;
			RECT 14.52 3.14 15 10.6 ;
			RECT 14.2 9.92 15 10.6 ;
			RECT 16.52 3.26 17.16 3.9 ;
			RECT 16.52 3.42 18.2 3.9 ;
			RECT 17.56 3.42 18.2 4.26 ;
			RECT 17.56 3.42 18.04 9.78 ;
			RECT 17.56 8.12 18.2 9.78 ;
			RECT 18.32 2.26 19.2 2.9 ;
			RECT 18.56 6.56 19.2 7.2 ;
			RECT 18.72 2.26 19.2 11.22 ;
			RECT 18.72 10.58 19.58 11.22 ;
			RECT 19.72 1.98 21.12 2.62 ;
			RECT 19.72 7.26 20.92 7.9 ;
			RECT 19.72 1.98 20.2 10.06 ;
			RECT 19.72 9.58 21.22 10.06 ;
			RECT 20.58 9.58 21.22 11.22 ;
			RECT 20.72 3.9 21.92 6.54 ;
			RECT 21.44 3.9 21.92 9.06 ;
			RECT 20.72 8.42 21.92 9.06 ;
			RECT 22.12 2 22.92 2.64 ;
			RECT 22.44 4.92 24.26 6.56 ;
			RECT 22.44 2 22.92 11.02 ;
			RECT 22.04 10.38 22.92 11.02 ;

	END

END MUX41XL

MACRO MUX41
	CLASS CORE ;
	FOREIGN MUX41 0 0  ;
	ORIGIN 0 0 ;
	SIZE 25.92 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.749 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 4.14 6.8 9.2 ;
			RECT 5.96 4.14 6.8 4.78 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.749 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 4.14 8.24 9.2 ;
			RECT 7.4 4.14 8.24 4.78 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.749 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 11.92 2.84 12.56 9.34 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.749 LAYER MTL1  ;
	END D
	PIN S1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 13.32 8.7 14 9.34 ;
			RECT 13.36 4.96 14 9.34 ;
			RECT 13.36 3.2 13.92 9.34 ;
			RECT 13.28 3.2 13.92 4.84 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.189 LAYER MTL1  ;
	END S1
	PIN S2
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 15.52 9.58 16.88 11.22 ;
			RECT 16.24 4.14 16.88 11.22 ;
			RECT 15.96 3.14 16.6 4.84 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.224 LAYER MTL1  ;
	END S2
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 24.88 1.98 25.52 11.02 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 25.92 13.68 ;
			RECT 23.44 10.34 24.08 13.68 ;
			RECT 17.5 10.74 18.14 13.68 ;
			RECT 12.8 9.92 13.44 13.68 ;
			RECT 6.84 10.02 7.48 13.68 ;
			RECT 0.96 10.12 1.6 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 25.92 1.46 ;
			RECT 22.76 -0.48 23.4 2.66 ;
			RECT 15.48 -0.48 16.12 2.62 ;
			RECT 12.4 -0.48 13.04 2.32 ;
			RECT 6.32 -0.48 6.96 3.4 ;
			RECT 1.04 -0.48 1.68 2.38 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1.56 3.26 2.84 3.9 ;
			RECT 2.36 3.26 2.84 10.8 ;
			RECT 2.36 10.16 3.04 10.8 ;
			RECT 3.36 2.54 4.12 7.12 ;
			RECT 3.78 6.48 4.44 10.8 ;
			RECT 4.8 2.54 5.44 3.18 ;
			RECT 4.96 2.54 5.44 10.86 ;
			RECT 4.96 10.22 6.08 10.86 ;
			RECT 7.96 1.98 8.6 3.62 ;
			RECT 7.96 3.14 9.24 3.62 ;
			RECT 8.76 3.14 9.24 10.66 ;
			RECT 8.24 10.02 9.24 10.66 ;
			RECT 9.36 1.98 10.24 2.62 ;
			RECT 9.76 1.98 10.24 10.54 ;
			RECT 9.76 5.2 10.4 10.54 ;
			RECT 10.76 1.98 11.4 2.62 ;
			RECT 10.92 1.98 11.4 10.66 ;
			RECT 10.92 10.02 12.04 10.66 ;
			RECT 14.04 2.02 14.96 2.68 ;
			RECT 14.48 2.02 14.96 3.62 ;
			RECT 14.52 7.56 15.32 8.2 ;
			RECT 14.52 3.14 15 10.6 ;
			RECT 14.2 9.92 15 10.6 ;
			RECT 17.12 2.06 18.04 2.7 ;
			RECT 17.4 2.06 18.04 9.34 ;
			RECT 17.5 8.2 18.14 9.98 ;
			RECT 18.56 3.7 19.2 4.34 ;
			RECT 18.56 6.56 19.2 7.2 ;
			RECT 18.72 3.7 19.2 11.22 ;
			RECT 18.72 10.58 19.58 11.22 ;
			RECT 19.08 1.98 20.24 2.62 ;
			RECT 19.72 1.98 20.24 7.7 ;
			RECT 19.72 6.06 20.56 7.7 ;
			RECT 19.72 1.98 20.2 10.06 ;
			RECT 19.72 9.58 21.22 10.06 ;
			RECT 20.58 9.58 21.22 11.22 ;
			RECT 20.8 1.98 21.92 2.62 ;
			RECT 20.76 3.54 21.92 5.18 ;
			RECT 21.44 1.98 21.92 8.86 ;
			RECT 20.72 8.22 21.92 8.86 ;
			RECT 22.76 3.66 23.4 6.3 ;
			RECT 22.44 4.66 23.78 6.3 ;
			RECT 22.44 4.66 22.92 11.02 ;
			RECT 22.04 10.38 22.92 11.02 ;

	END

END MUX41

MACRO MUX21XL
	CLASS CORE ;
	FOREIGN MUX21XL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 8.64 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.008 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 5.78 5.36 7.42 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.008 LAYER MTL1  ;
	END B
	PIN SA
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 4.96 1.04 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.584 LAYER MTL1  ;
	END SA
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.24 9.02 6.8 9.5 ;
			RECT 6.16 2.32 6.8 9.5 ;
			RECT 5.14 2.32 6.8 3.64 ;
			RECT 4.24 9.02 4.88 10.66 ;

		END 

		ANTENNADIFFAREA 2.912 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 8.64 13.68 ;
			RECT 6.64 10.02 7.28 13.68 ;
			RECT 1.84 9.76 2.48 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 8.64 1.46 ;
			RECT 7.56 -0.48 8.2 3.34 ;
			RECT 2.76 -0.48 3.4 3.34 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.76 1.98 1.76 2.62 ;
			RECT 1.12 1.98 1.76 4.34 ;
			RECT 1.12 3.86 3.48 4.34 ;
			RECT 3 3.86 3.48 8.28 ;
			RECT 1.36 7.64 3.48 8.28 ;
			RECT 1.36 7.64 1.86 9.24 ;
			RECT 0.4 8.76 1.86 9.24 ;
			RECT 0.4 8.76 1.04 10.3 ;

	END

END MUX21XL

MACRO MUX21
	CLASS CORE ;
	FOREIGN MUX21 0 0  ;
	ORIGIN 0 0 ;
	SIZE 11.52 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 5.28 5.36 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.261 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 5.28 8.24 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.261 LAYER MTL1  ;
	END B
	PIN SA
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 8.96 3.96 9.6 5.6 ;
			RECT 3.32 3.96 9.6 4.44 ;
			RECT 3.32 3.96 3.96 5.24 ;
			RECT 0.4 3.96 1.04 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 3.154 LAYER MTL1  ;
	END SA
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.24 8.24 11.12 8.94 ;
			RECT 10.48 2.96 11.12 8.94 ;
			RECT 5.2 2.96 11.12 3.44 ;
			RECT 5.64 8.24 6.28 10.94 ;
			RECT 5.2 2.8 5.84 3.44 ;

		END 

		ANTENNADIFFAREA 7.891 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 11.52 13.68 ;
			RECT 8.08 10.7 10.12 13.68 ;
			RECT 9.48 9.46 10.12 13.68 ;
			RECT 1.8 10.7 3.88 13.68 ;
			RECT 1.8 9.9 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 11.52 1.46 ;
			RECT 7.72 -0.48 8.36 2.44 ;
			RECT 2.8 -0.48 3.44 3.18 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.36 2.04 2.04 2.68 ;
			RECT 1.36 2.04 2.04 3.18 ;
			RECT 1.56 5.96 3 7.6 ;
			RECT 1.56 2.04 2.04 9.24 ;
			RECT 0.4 8.76 2.04 9.24 ;
			RECT 0.4 8.76 1.04 10.88 ;

	END

END MUX21

MACRO INVXL
	CLASS CORE ;
	FOREIGN INVXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 2.88 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 5.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.576 LAYER MTL1  ;
	END A
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 3.26 1.2 3.9 ;
			RECT 0.4 3.26 1.04 11.22 ;

		END 

		ANTENNADIFFAREA 1.614 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 2.88 13.68 ;
			RECT 1.8 10.58 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 2.88 1.46 ;
			RECT 0.56 -0.48 1.2 2.26 ;

		END 

	END gndd!

END INVXL

MACRO INV5
	CLASS CORE ;
	FOREIGN INV5 0 0  ;
	ORIGIN 0 0 ;
	SIZE 10.08 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 3.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 10.138 LAYER MTL1  ;
	END A
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.4 8.44 8.04 11.22 ;
			RECT 0.4 8.44 8.04 8.92 ;
			RECT 0.4 4.28 5.6 4.76 ;
			RECT 4.96 1.98 5.6 4.76 ;
			RECT 4.6 8.44 5.24 11.22 ;
			RECT 2.16 1.98 2.8 4.76 ;
			RECT 1.8 8.44 2.44 11.22 ;
			RECT 0.4 4.28 1.04 8.92 ;

		END 

		ANTENNADIFFAREA 14.643 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 10.08 13.68 ;
			RECT 8.8 8.44 9.44 13.68 ;
			RECT 6 9.44 6.64 13.68 ;
			RECT 3.2 9.44 3.84 13.68 ;
			RECT 0.4 9.44 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 10.08 1.46 ;
			RECT 6.36 -0.48 7 3.74 ;
			RECT 3.56 -0.48 4.2 3.76 ;
			RECT 0.76 -0.48 1.4 3.76 ;

		END 

	END gndd!

END INV5

MACRO INV4
	CLASS CORE ;
	FOREIGN INV4 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 3.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 6.84 LAYER MTL1  ;
	END A
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.6 8.44 5.24 11.22 ;
			RECT 0.4 8.44 5.24 8.92 ;
			RECT 0.4 4.28 2.8 4.76 ;
			RECT 2.16 1.98 2.8 4.76 ;
			RECT 1.8 8.44 2.44 11.22 ;
			RECT 0.4 4.28 1.04 8.92 ;

		END 

		ANTENNADIFFAREA 9.309 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 6 8.76 6.64 13.68 ;
			RECT 3.2 9.56 3.84 13.68 ;
			RECT 0.4 9.56 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 3.56 -0.48 4.2 3.44 ;
			RECT 0.76 -0.48 1.4 3.76 ;

		END 

	END gndd!

END INV4

MACRO INV3
	CLASS CORE ;
	FOREIGN INV3 0 0  ;
	ORIGIN 0 0 ;
	SIZE 5.76 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 3.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 5.069 LAYER MTL1  ;
	END A
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.6 8.7 5.24 11.22 ;
			RECT 0.4 8.7 5.24 9.18 ;
			RECT 0.4 3.82 2.8 4.3 ;
			RECT 2.16 1.98 2.8 4.3 ;
			RECT 1.8 8.7 2.44 11.22 ;
			RECT 0.4 3.82 1.04 9.18 ;

		END 

		ANTENNADIFFAREA 8.474 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 5.76 13.68 ;
			RECT 3.2 9.7 3.84 13.68 ;
			RECT 0.4 9.7 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 5.76 1.46 ;
			RECT 3.56 -0.48 4.2 3.3 ;
			RECT 0.76 -0.48 1.4 3.3 ;

		END 

	END gndd!

END INV3

MACRO INV2
	CLASS CORE ;
	FOREIGN INV2 0 0  ;
	ORIGIN 0 0 ;
	SIZE 4.32 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 3.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.534 LAYER MTL1  ;
	END A
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.8 8.62 2.44 11.22 ;
			RECT 0.4 8.62 2.44 9.1 ;
			RECT 0.4 1.98 1.4 3.82 ;
			RECT 0.4 1.98 1.04 9.1 ;

		END 

		ANTENNADIFFAREA 4.467 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 4.32 13.68 ;
			RECT 3.2 9.62 3.84 13.68 ;
			RECT 0.4 9.62 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 4.32 1.46 ;
			RECT 2.16 -0.48 2.8 3.3 ;

		END 

	END gndd!

END INV2

MACRO INV
	CLASS CORE ;
	FOREIGN INV 0 0  ;
	ORIGIN 0 0 ;
	SIZE 2.88 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 5.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.267 LAYER MTL1  ;
	END A
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 1.98 1.04 11.22 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 2.88 13.68 ;
			RECT 1.8 9.24 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 2.88 1.46 ;
			RECT 1.8 -0.48 2.44 2.64 ;

		END 

	END gndd!

END INV

MACRO HOLD
	CLASS CORE ;
	FOREIGN HOLD 0 0  ;
	ORIGIN 0 0 ;
	SIZE 4.32 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN O
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 2.36 7.68 3.92 9.54 ;
			RECT 3.28 3.06 3.92 9.54 ;
			RECT 3.12 3.06 3.92 3.7 ;
			RECT 1.32 7.68 3.92 8.34 ;

		END 

		ANTENNADIFFAREA 1.334 LAYER MTL1  ;
		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.461 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 4.32 13.68 ;
			RECT 2.4 10.58 3.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 4.32 1.46 ;
			RECT 0.72 -0.48 1.36 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.32 3.26 1.12 3.9 ;
			RECT 0.32 5.26 2.76 6.9 ;
			RECT 0.32 3.26 0.8 11.22 ;
			RECT 0.32 10.58 1.04 11.22 ;

	END

END HOLD

MACRO HADD
	CLASS CORE ;
	FOREIGN HADD 0 0  ;
	ORIGIN 0 0 ;
	SIZE 12.96 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.84 4.96 2.48 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.613 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.28 4.92 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.613 LAYER MTL1  ;
	END B
	PIN S
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 11.92 1.98 12.56 11.22 ;

		END 

		ANTENNADIFFAREA 3.232 LAYER MTL1  ;
	END S
	PIN C
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 9.04 3.54 10.2 4.18 ;
			RECT 9.04 9.02 9.76 11.22 ;
			RECT 9.04 3.54 9.68 11.22 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END C
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 12.96 13.68 ;
			RECT 10.52 9.02 11.16 13.68 ;
			RECT 7.68 10.7 8.32 13.68 ;
			RECT 3.84 9.9 4.48 13.68 ;
			RECT 1 9.9 1.64 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 12.96 1.46 ;
			RECT 9.16 -0.48 11.04 2.26 ;
			RECT 5.44 3.5 7.1 4.14 ;
			RECT 6.62 -0.48 7.1 4.14 ;
			RECT 0.72 -0.48 1.36 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1.88 1.98 6.04 2.62 ;
			RECT 1.88 1.98 2.38 3.26 ;
			RECT 0.68 2.78 2.38 3.26 ;
			RECT 0.68 2.78 1.32 3.98 ;
			RECT 3.16 3.22 4.92 3.86 ;
			RECT 4.44 3.22 4.92 5.14 ;
			RECT 4.44 4.66 7.16 5.14 ;
			RECT 5.68 8.7 7.16 9.18 ;
			RECT 6.52 4.66 7.16 9.18 ;
			RECT 2.4 8.9 6.16 9.38 ;
			RECT 2.4 8.9 3.04 10.54 ;
			RECT 7.72 1.98 8.36 2.62 ;
			RECT 7.88 4.98 8.52 6.62 ;
			RECT 7.88 1.98 8.36 10.18 ;
			RECT 6.68 9.7 8.36 10.18 ;
			RECT 6.68 9.7 7.16 11.22 ;
			RECT 6.28 10.58 7.16 11.22 ;

	END

END HADD

MACRO GNDTIE
	CLASS CORE ;
	FOREIGN GNDTIE 0 0  ;
	ORIGIN 0 0 ;
	SIZE 2.88 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 1.98 1.04 4.28 ;

		END 

		ANTENNADIFFAREA 0.986 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 2.88 13.68 ;
			RECT 1.7 10.94 2.36 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 2.88 1.46 ;
			RECT 1.8 -0.48 2.44 2.7 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.72 8.3 1.36 9.94 ;
			RECT 0.72 9.3 2.36 9.94 ;

	END

END GNDTIE

MACRO FSTDN8
	CLASS CORE SPACER ;
	FOREIGN FSTDN8 0 0  ;
	ORIGIN 0 0 ;
	SIZE 11.52 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 11.52 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 11.52 1.46 ;

		END 

	END gndd!

END FSTDN8

MACRO FSTDN4
	CLASS CORE SPACER ;
	FOREIGN FSTDN4 0 0  ;
	ORIGIN 0 0 ;
	SIZE 5.76 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 5.76 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 5.76 1.46 ;

		END 

	END gndd!

END FSTDN4

MACRO FSTDN2
	CLASS CORE SPACER ;
	FOREIGN FSTDN2 0 0  ;
	ORIGIN 0 0 ;
	SIZE 2.88 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 2.88 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 2.88 1.46 ;

		END 

	END gndd!

END FSTDN2

MACRO FSTDN16
	CLASS CORE SPACER ;
	FOREIGN FSTDN16 0 0  ;
	ORIGIN 0 0 ;
	SIZE 23.04 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 23.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 23.04 1.46 ;

		END 

	END gndd!

END FSTDN16

MACRO FSTDN
	CLASS CORE SPACER ;
	FOREIGN FSTDN 0 0  ;
	ORIGIN 0 0 ;
	SIZE 1.44 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 1.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 1.44 1.46 ;

		END 

	END gndd!

END FSTDN

MACRO FSTD8
	CLASS CORE SPACER ;
	FOREIGN FSTD8 0 0  ;
	ORIGIN 0 0 ;
	SIZE 11.52 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 11.52 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 11.52 1.46 ;

		END 

	END gndd!

END FSTD8

MACRO FSTD4
	CLASS CORE SPACER ;
	FOREIGN FSTD4 0 0  ;
	ORIGIN 0 0 ;
	SIZE 5.76 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 5.76 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 5.76 1.46 ;

		END 

	END gndd!

END FSTD4

MACRO FSTD2
	CLASS CORE SPACER ;
	FOREIGN FSTD2 0 0  ;
	ORIGIN 0 0 ;
	SIZE 2.88 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 2.88 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 2.88 1.46 ;

		END 

	END gndd!

END FSTD2

MACRO FSTD16
	CLASS CORE SPACER ;
	FOREIGN FSTD16 0 0  ;
	ORIGIN 0 0 ;
	SIZE 23.04 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 23.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 23.04 1.46 ;

		END 

	END gndd!

END FSTD16

MACRO FSTD
	CLASS CORE SPACER ;
	FOREIGN FSTD 0 0  ;
	ORIGIN 0 0 ;
	SIZE 1.44 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 1.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 1.44 1.46 ;

		END 

	END gndd!

END FSTD

MACRO FADD
	CLASS CORE ;
	FOREIGN FADD 0 0  ;
	ORIGIN 0 0 ;
	SIZE 28.8 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.28 4.92 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.837 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.84 4.96 2.48 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.837 LAYER MTL1  ;
	END B
	PIN CI
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 14.8 4.42 16.44 7.86 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.578 LAYER MTL1  ;
	END CI
	PIN S
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 27.76 2.32 28.4 11.22 ;
			RECT 26.24 2.96 28.4 3.64 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END S
	PIN CO
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 24.12 9 25.6 11.22 ;
			RECT 24.12 7.76 24.6 11.22 ;
			RECT 23.44 7.76 24.6 8.24 ;
			RECT 23.44 2.32 24.08 8.24 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END CO
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 28.8 13.68 ;
			RECT 26.36 9 27 13.68 ;
			RECT 22.94 8.76 23.6 13.68 ;
			RECT 19.1 8.38 19.74 13.68 ;
			RECT 17.38 10.78 18.04 13.68 ;
			RECT 11.32 8.5 11.96 13.68 ;
			RECT 5.64 9.86 6.28 13.68 ;
			RECT 2.8 9.76 3.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 28.8 1.46 ;
			RECT 24.84 -0.48 25.48 3.52 ;
			RECT 16.38 -0.48 17.02 2.62 ;
			RECT 12.54 -0.48 13.18 3.26 ;
			RECT 7.74 -0.48 8.38 3.26 ;
			RECT 3.7 -0.48 4.34 3.26 ;
			RECT 0.42 -0.48 1.12 3.12 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 4.24 8.86 7.72 9.34 ;
			RECT 4.24 8.86 4.88 10.54 ;
			RECT 7.08 8.86 7.72 10.54 ;
			RECT 2.06 2.62 2.7 4.26 ;
			RECT 2.06 3.78 5.58 4.26 ;
			RECT 5.1 3.78 5.58 5.42 ;
			RECT 5.1 4.78 8.62 5.42 ;
			RECT 7.32 4.78 7.96 8.3 ;
			RECT 3.24 7.66 7.96 8.3 ;
			RECT 3.24 7.66 3.72 9.24 ;
			RECT 0.4 8.76 3.72 9.24 ;
			RECT 0.4 8.76 1.04 10.58 ;
			RECT 6.1 2.62 6.74 4.26 ;
			RECT 6.1 3.78 9.62 4.26 ;
			RECT 9.14 3.78 9.62 6.9 ;
			RECT 8.48 6.18 12.66 6.9 ;
			RECT 8.48 6.18 9.12 10.54 ;
			RECT 9.92 7.42 12.96 7.9 ;
			RECT 12.48 7.42 12.96 11.22 ;
			RECT 9.92 7.42 10.56 10.38 ;
			RECT 12.48 9.38 13.36 11.22 ;
			RECT 15.6 9.38 16.24 11.22 ;
			RECT 12.48 10.74 16.24 11.22 ;
			RECT 10.14 2.62 10.78 4.78 ;
			RECT 10.14 4.3 13.96 4.78 ;
			RECT 16.96 4.5 19.48 5.14 ;
			RECT 13.48 4.3 13.96 8.86 ;
			RECT 16.96 4.5 17.44 8.86 ;
			RECT 13.48 8.38 17.44 8.86 ;
			RECT 14.2 8.38 14.84 9.88 ;
			RECT 14.94 2.62 15.58 3.62 ;
			RECT 14.94 3.14 20.48 3.62 ;
			RECT 19.84 3.14 20.48 3.78 ;
			RECT 20 3.14 20.48 7.86 ;
			RECT 18.1 7.22 20.48 7.86 ;
			RECT 18.1 7.22 18.58 10.02 ;
			RECT 17.56 9.38 18.58 10.02 ;
			RECT 20.36 1.98 22.08 2.62 ;
			RECT 21 1.98 22.08 3.62 ;
			RECT 21 1.98 21.48 9.2 ;
			RECT 20.56 8.56 21.48 9.2 ;

	END

END FADD

MACRO EXORXL
	CLASS CORE ;
	FOREIGN EXORXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 10.08 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 7.6 1.04 9.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.454 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 3.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.454 LAYER MTL1  ;
	END B
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 8.52 9.84 9.68 10.48 ;
			RECT 9.04 3.26 9.68 10.48 ;

		END 

		ANTENNADIFFAREA 1.701 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 10.08 13.68 ;
			RECT 7.08 9.66 7.72 13.68 ;
			RECT 3.2 9.86 3.84 13.68 ;
			RECT 0.4 9.86 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 10.08 1.46 ;
			RECT 8.92 -0.48 9.56 2.26 ;
			RECT 6.32 -0.48 6.96 2.26 ;
			RECT 3.04 -0.48 3.68 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 4.68 1.98 5.32 3.26 ;
			RECT 4.68 2.78 6.32 3.26 ;
			RECT 5.68 2.78 6.32 4.54 ;
			RECT 0.4 1.98 1.04 3.26 ;
			RECT 0.4 2.78 4.16 3.26 ;
			RECT 3.68 2.78 4.16 4.26 ;
			RECT 3.68 3.78 5.16 4.26 ;
			RECT 4.68 3.78 5.16 5.6 ;
			RECT 5.08 5.06 7.32 5.7 ;
			RECT 3.76 8.7 5.56 9.34 ;
			RECT 5.08 5.06 5.56 9.34 ;
			RECT 1.96 8.76 5.56 9.34 ;
			RECT 1.96 8.76 2.44 10.5 ;
			RECT 1.8 9.86 2.44 10.5 ;
			RECT 7.74 2.26 8.38 4.54 ;
			RECT 7.32 3.9 8.38 4.54 ;
			RECT 7.88 2.26 8.38 8.58 ;
			RECT 7.88 6.94 8.52 8.58 ;
			RECT 6.08 7.9 8.52 8.58 ;
			RECT 6.08 7.9 6.56 10.5 ;
			RECT 4.64 9.86 6.56 10.5 ;

	END

END EXORXL

MACRO EXOR
	CLASS CORE ;
	FOREIGN EXOR 0 0  ;
	ORIGIN 0 0 ;
	SIZE 10.08 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 7.58 1.04 9.22 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.598 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 5.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.598 LAYER MTL1  ;
	END B
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 9.04 1.98 9.68 8.9 ;
			RECT 8.52 8.26 9.16 10.12 ;
			RECT 8.88 1.98 9.68 2.62 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 10.08 13.68 ;
			RECT 7.08 8.9 7.72 13.68 ;
			RECT 3.2 9.76 3.84 13.68 ;
			RECT 0.4 9.76 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 10.08 1.46 ;
			RECT 7.28 -0.48 7.92 2.26 ;
			RECT 5.84 -0.48 6.48 2.62 ;
			RECT 3.04 -0.48 3.68 2.62 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 4.44 1.98 5.32 2.62 ;
			RECT 4.84 1.98 5.32 3.62 ;
			RECT 4.84 3.14 6.6 3.62 ;
			RECT 5.96 3.14 6.6 4.1 ;
			RECT 0.4 1.98 1.04 4.2 ;
			RECT 0.4 3.72 4.08 4.2 ;
			RECT 3.6 3.72 4.08 5.38 ;
			RECT 3.6 4.74 7.16 5.38 ;
			RECT 3.76 8.5 5.56 9.24 ;
			RECT 5.08 4.74 5.56 9.24 ;
			RECT 1.96 8.76 5.56 9.24 ;
			RECT 1.96 8.76 2.44 10.4 ;
			RECT 1.8 9.76 2.44 10.4 ;
			RECT 7.36 3.46 8.52 4.1 ;
			RECT 7.88 3.46 8.52 7.72 ;
			RECT 6.08 7.24 8.52 7.72 ;
			RECT 6.08 7.24 6.56 10.4 ;
			RECT 4.64 9.76 6.56 10.4 ;

	END

END EXOR

MACRO EXNORXL
	CLASS CORE ;
	FOREIGN EXNORXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 8.64 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 7.6 1.04 9.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.541 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 5.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.541 LAYER MTL1  ;
	END B
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.38 3.06 8.24 3.7 ;
			RECT 6.06 6.28 7.86 6.92 ;
			RECT 7.38 3.06 7.86 6.92 ;
			RECT 6.06 6.28 6.8 8.24 ;
			RECT 4.64 10.2 6.56 10.84 ;
			RECT 6.06 6.28 6.56 10.84 ;

		END 

		ANTENNADIFFAREA 2.536 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 8.64 13.68 ;
			RECT 7.08 10.08 7.72 13.68 ;
			RECT 3.2 10.2 3.84 13.68 ;
			RECT 0.4 10.08 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 8.64 1.46 ;
			RECT 6.08 -0.48 6.72 2.26 ;
			RECT 3.04 -0.48 3.68 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 1.98 1.04 3.26 ;
			RECT 0.4 2.78 4.04 3.26 ;
			RECT 3.56 4.62 6.32 5.26 ;
			RECT 3.56 2.78 4.04 9.68 ;
			RECT 3.56 8.04 4.32 9.68 ;
			RECT 1.8 9.04 4.32 9.68 ;
			RECT 1.8 9.04 2.44 10.72 ;
			RECT 4.56 1.98 5.2 3.26 ;
			RECT 4.56 2.78 6.86 3.26 ;
			RECT 6.2 2.78 6.86 3.7 ;

	END

END EXNORXL

MACRO EXNOR
	CLASS CORE ;
	FOREIGN EXNOR 0 0  ;
	ORIGIN 0 0 ;
	SIZE 12.96 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 7.46 1.04 9.1 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.995 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.96 3.48 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.995 LAYER MTL1  ;
	END B
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 5 4.96 10.48 5.6 ;
			RECT 9.84 1.98 10.48 5.6 ;
			RECT 4.64 10.74 8.12 11.22 ;
			RECT 7.48 9.8 8.12 11.22 ;
			RECT 4.64 8.6 5.48 11.22 ;
			RECT 5 4.96 5.48 11.22 ;

		END 

		ANTENNADIFFAREA 5.947 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 12.96 13.68 ;
			RECT 10.28 9.8 10.92 13.68 ;
			RECT 3.2 9.78 3.84 13.68 ;
			RECT 0.4 9.72 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 12.96 1.46 ;
			RECT 7 -0.48 7.64 2.26 ;
			RECT 4.16 -0.48 4.8 2.34 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 8.16 1.98 9.08 2.62 ;
			RECT 5.6 1.98 6.26 3.26 ;
			RECT 8.16 1.98 8.64 3.26 ;
			RECT 5.6 2.78 8.64 3.26 ;
			RECT 1.62 1.98 2.26 3.46 ;
			RECT 1.62 2.98 4.48 3.46 ;
			RECT 4 3.78 9.12 4.42 ;
			RECT 4 2.98 4.48 8.08 ;
			RECT 3.64 6.34 4.12 9.24 ;
			RECT 1.8 8.76 4.12 9.24 ;
			RECT 1.8 8.76 2.44 10.36 ;
			RECT 6.08 8.76 12.32 9.28 ;
			RECT 6.08 8.76 6.72 10.06 ;
			RECT 8.88 8.76 9.52 10.06 ;
			RECT 11.68 8.76 12.32 10.06 ;

	END

END EXNOR

MACRO DLLRL
	CLASS CORE ;
	FOREIGN DLLRL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 20.16 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 3.96 1.04 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.109 LAYER MTL1  ;
	END D
	PIN ENB
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 3.96 6.8 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.936 LAYER MTL1  ;
	END ENB
	PIN RB
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 2.48 7.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.037 LAYER MTL1  ;
	END RB
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 19.12 2.8 19.76 10.88 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END Q
	PIN QB
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 16.24 8.34 17 10.66 ;
			RECT 16.24 2.8 16.98 3.44 ;
			RECT 16.24 2.8 16.88 10.88 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END QB
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 20.16 13.68 ;
			RECT 17.72 8.34 18.36 13.68 ;
			RECT 13.44 10.7 14.08 13.68 ;
			RECT 7.72 10.74 8.36 13.68 ;
			RECT 4.44 10.7 5.08 13.68 ;
			RECT 0.4 9.7 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 20.16 1.46 ;
			RECT 17.72 -0.48 18.36 3.44 ;
			RECT 13.24 -0.48 13.88 3.06 ;
			RECT 6.64 -0.48 7.28 3.18 ;
			RECT 0.4 -0.48 1.04 3.36 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 4.96 2.54 5.88 3.18 ;
			RECT 4.96 2.54 5.44 4.4 ;
			RECT 4 3.92 5.44 4.4 ;
			RECT 4 3.92 4.64 9.18 ;
			RECT 8.2 7.74 8.84 9.18 ;
			RECT 4 8.54 8.84 9.18 ;
			RECT 8.16 2.54 9.08 3.18 ;
			RECT 8.58 2.54 9.08 4.18 ;
			RECT 8.58 3.7 10.44 4.18 ;
			RECT 9.36 3.7 10.44 5.34 ;
			RECT 5.44 6.38 9.84 6.86 ;
			RECT 5.44 6.38 6.08 8.02 ;
			RECT 9.36 3.7 9.84 9.18 ;
			RECT 9.36 8.54 10 9.18 ;
			RECT 9.6 2.54 11.44 3.18 ;
			RECT 3 2.7 4.44 3.34 ;
			RECT 3 2.7 3.48 10.18 ;
			RECT 2.8 9.7 11.44 10.18 ;
			RECT 2.8 9.58 3.44 11.22 ;
			RECT 10.96 2.54 11.44 11.22 ;
			RECT 9.8 9.7 11.44 11.22 ;
			RECT 14.88 2.42 15.52 4.06 ;
			RECT 12.6 3.58 15.52 4.06 ;
			RECT 12.6 3.58 13.24 10.18 ;
			RECT 12.6 9.7 15.48 10.18 ;
			RECT 14.84 9.7 15.48 11.22 ;

	END

END DLLRL

MACRO DLL
	CLASS CORE ;
	FOREIGN DLL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 18.72 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.08 LAYER MTL1  ;
	END D
	PIN ENB
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 3.16 6.8 9.56 ;
			RECT 5.44 7.96 6.8 8.92 ;
			RECT 5.44 3.16 6.8 3.8 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.936 LAYER MTL1  ;
	END ENB
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 16.94 10.58 18.32 11.22 ;
			RECT 17.68 2.08 18.32 11.22 ;
			RECT 17.48 2.08 18.32 2.72 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END Q
	PIN QB
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 14.14 9.22 16.88 9.7 ;
			RECT 16.24 3.14 16.88 9.7 ;
			RECT 14.68 3.14 16.88 3.62 ;
			RECT 14.68 1.98 15.32 3.62 ;
			RECT 14.14 9.22 14.78 11.22 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END QB
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 18.72 13.68 ;
			RECT 15.54 10.22 16.18 13.68 ;
			RECT 11.16 9.58 11.8 13.68 ;
			RECT 5.64 10.12 6.28 13.68 ;
			RECT 0.4 10.08 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 18.72 1.46 ;
			RECT 16.08 -0.48 16.72 2.62 ;
			RECT 11.6 -0.48 12.24 2.62 ;
			RECT 5.84 -0.48 6.48 2.54 ;
			RECT 0.4 -0.48 1.04 2.34 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 2.76 1.98 3.44 2.62 ;
			RECT 2.76 4.52 3.92 5.16 ;
			RECT 2.76 1.98 3.24 11.22 ;
			RECT 2.76 9.58 3.44 11.22 ;
			RECT 4.44 1.98 5.08 2.62 ;
			RECT 3.96 3.16 4.92 3.8 ;
			RECT 4.44 5.52 5.28 6.16 ;
			RECT 4.44 1.98 4.92 10.82 ;
			RECT 4.24 9.58 4.92 10.82 ;
			RECT 7.52 1.98 8.16 3.8 ;
			RECT 7.52 3.14 9.64 3.8 ;
			RECT 8.64 3.14 9.28 7.6 ;
			RECT 7.52 6.96 9.28 7.6 ;
			RECT 7.52 6.96 8.16 8.6 ;
			RECT 7.52 6.96 8 11.22 ;
			RECT 7.08 10.52 8 11.22 ;
			RECT 8.96 1.98 10.64 2.62 ;
			RECT 10 4.52 10.64 11.22 ;
			RECT 10.16 1.98 10.64 11.22 ;
			RECT 8.52 10.58 10.64 11.22 ;
			RECT 13.14 2.58 13.88 4.78 ;
			RECT 13.14 4.14 15.72 4.78 ;
			RECT 13.14 7.02 13.8 8.66 ;
			RECT 13.14 2.58 13.62 10.5 ;
			RECT 12.7 9.86 13.62 10.5 ;

	END

END DLL

MACRO DLHRL
	CLASS CORE ;
	FOREIGN DLHRL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 20.16 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 3.96 1.04 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.109 LAYER MTL1  ;
	END D
	PIN EN
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER MTL1 ;
			RECT 5.14 4.96 6.8 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.08 LAYER MTL1  ;
	END EN
	PIN RB
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 2.48 7.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.037 LAYER MTL1  ;
	END RB
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 19.12 2.8 19.76 10.88 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END Q
	PIN QB
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 16.24 8.34 17 10.66 ;
			RECT 16.24 2.8 16.98 3.44 ;
			RECT 16.24 2.8 16.88 10.88 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END QB
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 20.16 13.68 ;
			RECT 17.72 8.34 18.36 13.68 ;
			RECT 13.24 10.7 13.88 13.68 ;
			RECT 7.52 10.74 8.16 13.68 ;
			RECT 4.44 10.7 5.08 13.68 ;
			RECT 0.4 9.7 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 20.16 1.46 ;
			RECT 17.72 -0.48 18.36 3.44 ;
			RECT 13.24 -0.48 13.88 2.62 ;
			RECT 6.64 -0.48 7.28 3.18 ;
			RECT 0.4 -0.48 1.04 3.36 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 4.96 2.54 5.88 3.18 ;
			RECT 4.96 2.54 5.44 4.4 ;
			RECT 4 3.92 5.44 4.4 ;
			RECT 4 3.92 4.48 9.18 ;
			RECT 8 7.74 8.64 9.18 ;
			RECT 4 8.54 8.64 9.18 ;
			RECT 8.16 2.54 9.08 3.18 ;
			RECT 8.58 3.14 11.08 3.62 ;
			RECT 5 6.74 11.08 7.22 ;
			RECT 5 6.74 5.64 7.38 ;
			RECT 10.58 3.14 11.08 9.18 ;
			RECT 9.16 6.74 11.08 9.18 ;
			RECT 9.6 1.98 12.08 2.62 ;
			RECT 3 2.7 4.44 3.34 ;
			RECT 3 2.7 3.48 10.18 ;
			RECT 2.8 9.7 12.08 10.18 ;
			RECT 11.6 1.98 12.08 10.86 ;
			RECT 9.6 9.7 12.08 10.86 ;
			RECT 2.8 9.58 3.44 11.22 ;
			RECT 9.6 9.7 10.24 11.22 ;
			RECT 14.88 2.42 15.52 3.62 ;
			RECT 12.6 3.14 15.52 3.62 ;
			RECT 12.6 3.14 13.24 10.18 ;
			RECT 12.6 9.7 15.28 10.18 ;
			RECT 14.64 9.7 15.28 11.22 ;

	END

END DLHRL

MACRO DLH
	CLASS CORE ;
	FOREIGN DLH 0 0  ;
	ORIGIN 0 0 ;
	SIZE 18.72 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.08 LAYER MTL1  ;
	END D
	PIN EN
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER MTL1 ;
			RECT 5.44 8.24 7.08 8.92 ;
			RECT 5.44 8.24 6.8 9.56 ;
			RECT 6.16 3.16 6.8 9.56 ;
			RECT 5.44 3.16 6.8 4.96 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.08 LAYER MTL1  ;
	END EN
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 16.94 10.58 18.32 11.22 ;
			RECT 17.68 2.08 18.32 11.22 ;
			RECT 17.48 2.08 18.32 2.72 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END Q
	PIN QB
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 14.14 9.22 16.88 9.7 ;
			RECT 16.24 3.14 16.88 9.7 ;
			RECT 14.68 3.14 16.88 3.62 ;
			RECT 14.68 1.98 15.32 3.62 ;
			RECT 14.14 9.22 14.78 11.22 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END QB
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 18.72 13.68 ;
			RECT 15.54 10.22 16.18 13.68 ;
			RECT 11.16 9.58 11.8 13.68 ;
			RECT 5.64 10.12 6.28 13.68 ;
			RECT 0.4 10.08 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 18.72 1.46 ;
			RECT 16.08 -0.48 16.72 2.62 ;
			RECT 11.6 -0.48 12.24 2.62 ;
			RECT 5.84 -0.48 6.48 2.52 ;
			RECT 0.4 -0.48 1.04 2.34 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 2.76 1.98 3.44 2.62 ;
			RECT 2.76 5.56 3.92 6.2 ;
			RECT 2.76 1.98 3.24 11.22 ;
			RECT 2.76 9.58 3.44 11.22 ;
			RECT 4.44 1.98 5.08 2.62 ;
			RECT 3.96 3.16 4.92 4.8 ;
			RECT 3.76 8.42 4.92 9.06 ;
			RECT 4.44 1.98 4.92 11.22 ;
			RECT 4.24 8.42 4.92 11.22 ;
			RECT 7.52 2.16 8.16 3.72 ;
			RECT 7.52 3.14 9.28 3.72 ;
			RECT 8.64 3.14 9.28 10.06 ;
			RECT 7.52 9.58 9.28 10.06 ;
			RECT 7.52 9.58 8 11.22 ;
			RECT 7.08 10.52 8 11.22 ;
			RECT 8.96 1.98 10.64 2.62 ;
			RECT 10 1.98 10.64 11.22 ;
			RECT 8.52 10.58 10.64 11.22 ;
			RECT 13.14 2.58 13.88 4.78 ;
			RECT 13.14 4.14 15.72 4.78 ;
			RECT 13.14 7.02 13.8 8.66 ;
			RECT 13.14 2.58 13.62 10.5 ;
			RECT 12.7 9.86 13.62 10.5 ;

	END

END DLH

MACRO DFSSLQ
	CLASS CORE ;
	FOREIGN DFSSLQ 0 0  ;
	ORIGIN 0 0 ;
	SIZE 28.8 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN C
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER MTL1 ;
			RECT 18.2 6.28 18.84 9.04 ;
			RECT 16.24 6.28 18.84 6.92 ;
			RECT 16.24 4.96 17.64 6.92 ;
			RECT 17 3.54 17.64 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.821 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 3.96 1.04 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.662 LAYER MTL1  ;
	END D
	PIN SB
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 8.76 9.22 10.4 9.86 ;
			RECT 9.04 3.14 9.76 4.78 ;
			RECT 9.04 3.14 9.68 9.86 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.57 LAYER MTL1  ;
	END SB
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 27.76 1.98 28.4 11.22 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END Q
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 28.8 13.68 ;
			RECT 26.36 9.12 27 13.68 ;
			RECT 24.92 10.58 25.56 13.68 ;
			RECT 19.12 10.68 19.76 13.68 ;
			RECT 13.84 10.32 14.48 13.68 ;
			RECT 10.76 10.58 11.4 13.68 ;
			RECT 8.16 10.58 8.8 13.68 ;
			RECT 5.36 10.7 6 13.68 ;
			RECT 0.4 10.7 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 28.8 1.46 ;
			RECT 26.36 -0.48 27 2.5 ;
			RECT 20.82 -0.48 21.46 1.8 ;
			RECT 16 -0.48 16.64 2.54 ;
			RECT 9.76 -0.48 10.4 2.62 ;
			RECT 5.68 -0.48 6.32 2.62 ;
			RECT 0.4 -0.48 1.04 2.62 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 2.56 3.14 4.04 4.78 ;
			RECT 2.56 3.14 3.04 9.18 ;
			RECT 2.36 8.54 3.04 9.18 ;
			RECT 1.56 1.98 3.68 2.62 ;
			RECT 4.6 3.14 6.68 3.8 ;
			RECT 1.56 1.98 2.04 8.02 ;
			RECT 1.36 7.54 1.84 10.18 ;
			RECT 4.6 9.22 6.36 9.86 ;
			RECT 4.6 3.14 5.08 10.18 ;
			RECT 1.36 9.7 5.08 10.18 ;
			RECT 2.8 9.7 3.44 11.22 ;
			RECT 7.12 1.98 7.76 2.62 ;
			RECT 7.2 1.98 7.68 5 ;
			RECT 5.6 4.52 7.36 5.16 ;
			RECT 5.6 4.52 6.08 8.5 ;
			RECT 5.6 7.86 7.52 8.5 ;
			RECT 6.88 7.86 7.52 11.22 ;
			RECT 6.76 10.58 7.52 11.22 ;
			RECT 10.92 1.98 12.8 2.62 ;
			RECT 10.92 1.98 11.4 6.18 ;
			RECT 10.92 5.54 12.84 6.18 ;
			RECT 11.92 5.54 12.4 10.7 ;
			RECT 11.92 10.06 13.04 10.7 ;
			RECT 14.36 3.54 16.14 4.18 ;
			RECT 14.36 3.54 14.84 8.54 ;
			RECT 14.36 7.9 15 8.54 ;
			RECT 13.36 1.98 14.24 2.62 ;
			RECT 11.92 3.52 13.84 4.16 ;
			RECT 16.24 8.26 17.4 8.9 ;
			RECT 13.36 1.98 13.84 9.54 ;
			RECT 12.92 8.9 13.84 9.54 ;
			RECT 12.92 9.06 16.88 9.54 ;
			RECT 16.24 8.26 16.88 11.22 ;
			RECT 17.52 1.98 18.66 2.62 ;
			RECT 18.18 1.98 18.66 3.96 ;
			RECT 18.18 3.32 19.88 3.96 ;
			RECT 19.4 8.4 20.32 9.06 ;
			RECT 19.4 3.32 19.88 10.04 ;
			RECT 17.68 9.56 19.88 10.04 ;
			RECT 17.68 9.56 18.36 11.22 ;
			RECT 19.18 1.98 19.82 2.8 ;
			RECT 19.18 2.32 21.82 2.8 ;
			RECT 20.48 4.54 21.82 5.18 ;
			RECT 21.34 2.32 21.82 10.06 ;
			RECT 21.34 9.42 23.24 10.06 ;
			RECT 20.96 9.58 21.44 11.22 ;
			RECT 20.52 10.58 21.44 11.22 ;
			RECT 23.48 1.98 24.36 2.62 ;
			RECT 22.34 7.06 24.36 8.7 ;
			RECT 23.88 1.98 24.36 11.22 ;
			RECT 21.96 10.58 24.36 11.22 ;
			RECT 24.92 3.66 26.16 4.3 ;
			RECT 24.92 6.18 25.64 7.82 ;
			RECT 24.92 3.66 25.56 9.74 ;

	END

END DFSSLQ

MACRO DFSRLSLQ
	CLASS CORE ;
	FOREIGN DFSRLSLQ 0 0  ;
	ORIGIN 0 0 ;
	SIZE 34.56 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN C
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER MTL1 ;
			RECT 23.96 6.28 24.6 9.04 ;
			RECT 22 7.6 24.6 8.24 ;
			RECT 22.42 6.28 24.6 8.24 ;
			RECT 22.42 3.76 23.06 8.24 ;
			RECT 22 6.28 24.6 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.821 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.662 LAYER MTL1  ;
	END D
	PIN RB
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 12.08 4.54 12.76 5.18 ;
			RECT 11.14 6.28 12.56 8.24 ;
			RECT 12.08 4.54 12.56 8.24 ;
			RECT 11.14 6.28 11.96 9.56 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.562 LAYER MTL1  ;
	END RB
	PIN SB
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 14.32 8.9 16 9.54 ;
			RECT 15.52 5.54 16 9.54 ;
			RECT 14.28 5.54 16 6.18 ;
			RECT 4.6 3.14 6.68 3.8 ;
			RECT 4.6 9.46 6.36 10.14 ;
			RECT 4.6 7.6 5.36 10.14 ;
			RECT 4.6 6.28 5.36 6.92 ;
			RECT 4.6 3.14 5.08 10.14 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.872 LAYER MTL1  ;
	END SB
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 33.52 1.98 34.16 11.22 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END Q
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 34.56 13.68 ;
			RECT 32.12 9.26 32.76 13.68 ;
			RECT 30.68 10.58 31.32 13.68 ;
			RECT 24.88 10.68 25.52 13.68 ;
			RECT 19.6 10.32 20.24 13.68 ;
			RECT 15.24 11.06 15.88 13.68 ;
			RECT 10.32 10.58 10.96 13.68 ;
			RECT 5.36 11.66 6 13.68 ;
			RECT 0.4 10.7 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 34.56 1.46 ;
			RECT 32.12 -0.48 32.76 2.66 ;
			RECT 26.58 -0.48 27.22 1.8 ;
			RECT 21.56 -0.48 22.2 2.54 ;
			RECT 13.4 -0.48 14.04 2.5 ;
			RECT 5.68 -0.48 6.32 2.58 ;
			RECT 0.4 -0.48 1.04 2.62 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 2.56 3.14 4.04 4.78 ;
			RECT 2.56 3.14 3.04 9.18 ;
			RECT 2.36 8.54 3.04 9.18 ;
			RECT 8.6 2.98 9.24 5 ;
			RECT 5.6 4.52 9.24 5 ;
			RECT 5.6 4.52 7.56 5.16 ;
			RECT 7.08 4.52 7.56 8.54 ;
			RECT 7.28 7.9 7.92 10.14 ;
			RECT 1.56 1.98 3.68 2.62 ;
			RECT 9.76 3.14 10.4 3.78 ;
			RECT 1.56 1.98 2.04 8.02 ;
			RECT 9.76 3.14 10.24 9.7 ;
			RECT 8.44 9.06 10.24 9.7 ;
			RECT 1.36 7.54 1.84 10.18 ;
			RECT 1.56 9.7 2.04 11.22 ;
			RECT 8.44 9.06 8.92 11.14 ;
			RECT 1.56 10.66 8.92 11.14 ;
			RECT 1.56 10.58 3.44 11.22 ;
			RECT 7.08 1.98 10.76 2.46 ;
			RECT 7.08 1.98 7.72 2.62 ;
			RECT 10.12 1.98 10.76 2.62 ;
			RECT 11.76 1.98 12.4 4.02 ;
			RECT 10.92 3.54 15.8 4.02 ;
			RECT 15.32 3.54 15.8 4.78 ;
			RECT 15.32 4.14 15.96 4.78 ;
			RECT 10.92 3.54 11.4 5.18 ;
			RECT 10.76 4.54 11.4 5.18 ;
			RECT 13.28 3.54 13.76 9.54 ;
			RECT 12.48 8.9 13.76 9.54 ;
			RECT 12.48 8.9 13 11.22 ;
			RECT 11.88 10.58 13 11.22 ;
			RECT 16.32 2.98 17 3.62 ;
			RECT 16.52 5.54 18.28 6.18 ;
			RECT 16.52 2.98 17 10.54 ;
			RECT 13.72 10.06 18.28 10.54 ;
			RECT 13.72 10.06 14.36 11.22 ;
			RECT 17.64 10.06 18.28 11.22 ;
			RECT 14.8 1.98 18.36 2.46 ;
			RECT 14.8 1.98 15.44 2.62 ;
			RECT 17.72 1.98 18.36 3.34 ;
			RECT 20 3.76 21.7 4.4 ;
			RECT 20 3.76 20.48 8.54 ;
			RECT 20 7.9 20.64 8.54 ;
			RECT 19 1.98 19.8 2.62 ;
			RECT 17.52 4.18 19.48 4.82 ;
			RECT 19 1.98 19.48 9.54 ;
			RECT 18.64 8.9 19.48 9.54 ;
			RECT 22.04 8.9 23.16 9.54 ;
			RECT 18.64 9.06 23.16 9.54 ;
			RECT 22 9.06 22.64 11.22 ;
			RECT 23.2 1.98 24.06 2.62 ;
			RECT 23.58 1.98 24.06 4.62 ;
			RECT 23.58 4.14 26.58 4.62 ;
			RECT 25.94 3.36 26.58 5 ;
			RECT 25.56 8.4 26.4 9.06 ;
			RECT 25.56 4.14 26.04 10.04 ;
			RECT 23.68 9.56 26.04 10.04 ;
			RECT 23.68 9.56 24.16 11.22 ;
			RECT 23.44 10.5 24.16 11.22 ;
			RECT 24.58 1.98 25.58 2.8 ;
			RECT 24.58 2.32 27.58 2.8 ;
			RECT 24.58 1.98 25.22 3.62 ;
			RECT 27.1 2.32 27.58 10.06 ;
			RECT 27.1 9.42 29 10.06 ;
			RECT 26.72 9.58 27.2 11.22 ;
			RECT 26.28 10.58 27.2 11.22 ;
			RECT 28.1 1.98 29.88 2.62 ;
			RECT 28.1 1.98 28.74 8.9 ;
			RECT 28.1 8.42 30 8.9 ;
			RECT 29.52 8.42 30 11.22 ;
			RECT 27.72 10.58 30 11.22 ;
			RECT 29.26 3.66 31.92 4.3 ;
			RECT 29.26 3.66 29.74 7.5 ;
			RECT 29.26 7.02 31.36 7.5 ;
			RECT 30.64 7.02 31.36 9.74 ;

	END

END DFSRLSLQ

MACRO DFSRLQ
	CLASS CORE ;
	FOREIGN DFSRLQ 0 0  ;
	ORIGIN 0 0 ;
	SIZE 33.12 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN C
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER MTL1 ;
			RECT 22.52 6.28 23.16 9.04 ;
			RECT 20.56 7.6 23.16 8.24 ;
			RECT 20.98 6.28 23.16 8.24 ;
			RECT 20.98 3.76 21.62 8.24 ;
			RECT 20.56 6.28 23.16 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.821 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 5.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.691 LAYER MTL1  ;
	END D
	PIN RB
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 12.36 8.9 14 9.56 ;
			RECT 13.36 3.14 14 9.56 ;
			RECT 12.84 3.14 14 4.78 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.562 LAYER MTL1  ;
	END RB
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 32.08 1.98 32.72 11.22 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END Q
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 33.12 13.68 ;
			RECT 30.68 9.1 31.32 13.68 ;
			RECT 29.24 10.58 29.88 13.68 ;
			RECT 23.44 10.68 24.08 13.68 ;
			RECT 18.16 10.74 18.8 13.68 ;
			RECT 13.6 10.38 14.24 13.68 ;
			RECT 9.64 11.22 10.28 13.68 ;
			RECT 5.8 10.7 6.44 13.68 ;
			RECT 0.96 10.7 1.6 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 33.12 1.46 ;
			RECT 30.68 -0.48 31.32 2.66 ;
			RECT 25.14 -0.48 25.78 1.8 ;
			RECT 20.12 -0.48 20.76 2.82 ;
			RECT 16.26 -0.48 16.92 2.62 ;
			RECT 13.48 -0.48 14.12 2.62 ;
			RECT 10.4 -0.48 11.04 2.14 ;
			RECT 7.12 -0.48 7.76 1.78 ;
			RECT 1.82 -0.48 2.46 2.3 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 5.08 3.3 5.72 9.18 ;
			RECT 2.92 8.54 5.72 9.18 ;
			RECT 8.76 1.98 9.4 2.78 ;
			RECT 7.4 2.3 9.4 2.78 ;
			RECT 7.4 2.3 8.04 8.34 ;
			RECT 9.56 7.7 10.2 10.7 ;
			RECT 7.24 10.22 10.2 10.7 ;
			RECT 7.24 10.22 7.94 10.86 ;
			RECT 4.46 1.98 5.14 2.78 ;
			RECT 4.46 2.3 6.72 2.78 ;
			RECT 9.92 2.66 10.56 3.78 ;
			RECT 8.56 3.3 10.56 3.78 ;
			RECT 6.24 9.06 9.04 9.7 ;
			RECT 8.56 3.3 9.04 9.7 ;
			RECT 6.24 2.3 6.72 10.18 ;
			RECT 3.36 9.7 6.72 10.18 ;
			RECT 3.36 9.7 4 11.22 ;
			RECT 11.56 1.98 12.48 2.62 ;
			RECT 11.56 1.98 12.04 4.94 ;
			RECT 9.72 4.3 12.04 4.94 ;
			RECT 10.72 4.3 11.2 10.7 ;
			RECT 11.16 10.22 12.8 11.22 ;
			RECT 14.88 1.98 15.74 2.62 ;
			RECT 15.26 1.98 15.74 3.62 ;
			RECT 15.7 3.14 16.52 5.62 ;
			RECT 16 3.14 16.52 11.22 ;
			RECT 16 9.44 16.64 11.22 ;
			RECT 18.44 3.76 20.26 4.4 ;
			RECT 18.44 3.76 18.92 8.38 ;
			RECT 18.2 7.7 18.92 8.38 ;
			RECT 17.44 1.98 18.36 2.62 ;
			RECT 17.44 1.98 17.92 4.38 ;
			RECT 20.56 8.9 21.72 9.54 ;
			RECT 17.2 3.74 17.68 10.22 ;
			RECT 17.2 9.56 21.2 10.22 ;
			RECT 20.56 8.9 21.2 11.22 ;
			RECT 21.76 1.98 22.62 2.62 ;
			RECT 22.14 1.98 22.62 4.62 ;
			RECT 24.5 3.36 25.14 4.62 ;
			RECT 22.14 4.14 25.14 4.62 ;
			RECT 24.16 7.42 24.96 9.06 ;
			RECT 24.16 4.14 24.64 10.04 ;
			RECT 22.24 9.56 24.64 10.04 ;
			RECT 22.24 9.56 22.72 11.22 ;
			RECT 22 10.5 22.72 11.22 ;
			RECT 23.14 1.98 24.14 2.8 ;
			RECT 23.14 2.32 26.14 2.8 ;
			RECT 23.14 1.98 23.78 3.62 ;
			RECT 25.66 2.32 26.14 10.06 ;
			RECT 25.66 8.9 26.36 10.06 ;
			RECT 25.28 9.58 25.76 11.22 ;
			RECT 24.84 10.58 25.76 11.22 ;
			RECT 26.88 1.98 28.44 2.62 ;
			RECT 26.66 6.52 27.36 8.16 ;
			RECT 26.88 1.98 27.36 11.22 ;
			RECT 26.28 10.58 27.36 11.22 ;
			RECT 27.88 3.66 30.48 4.3 ;
			RECT 27.88 3.66 28.36 7.5 ;
			RECT 27.88 7.02 29.92 7.5 ;
			RECT 29.14 7.02 29.92 9.74 ;

	END

END DFSRLQ

MACRO DFSQ
	CLASS CORE ;
	FOREIGN DFSQ 0 0  ;
	ORIGIN 0 0 ;
	SIZE 25.92 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN C
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER MTL1 ;
			RECT 14.8 7.6 16.88 8.24 ;
			RECT 15.22 6.28 16.88 8.24 ;
			RECT 16.04 6.28 16.68 9.04 ;
			RECT 15.22 3.76 15.86 8.24 ;
			RECT 14.8 6.28 16.88 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.821 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 6.28 1.04 7.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.648 LAYER MTL1  ;
	END D
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 24.88 1.98 25.52 11.22 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END Q
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 25.92 13.68 ;
			RECT 22.08 10.58 24.12 13.68 ;
			RECT 23.48 9.1 24.12 13.68 ;
			RECT 16.6 10.68 17.24 13.68 ;
			RECT 11.32 10.14 11.96 13.68 ;
			RECT 8.28 10.38 8.92 13.68 ;
			RECT 5.24 10.7 5.88 13.68 ;
			RECT 0.4 10.7 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 25.92 1.46 ;
			RECT 23.48 -0.48 24.12 2.26 ;
			RECT 19.38 -0.48 20.02 1.8 ;
			RECT 14.36 -0.48 15 2.82 ;
			RECT 8.86 -0.48 9.5 2.14 ;
			RECT 5.78 -0.48 6.42 1.78 ;
			RECT 0.48 -0.48 1.12 2.3 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 3.48 3.3 4.12 8.9 ;
			RECT 2.36 8.22 4.12 8.9 ;
			RECT 2.36 8.22 3 9.86 ;
			RECT 3.12 1.98 3.8 2.78 ;
			RECT 3.12 2.3 5.22 2.78 ;
			RECT 4.74 4.04 5.78 5.72 ;
			RECT 4.74 2.3 5.22 10.18 ;
			RECT 4.04 9.7 5.22 10.18 ;
			RECT 4.04 9.7 4.52 11.22 ;
			RECT 2.8 10.58 4.52 11.22 ;
			RECT 7.22 1.98 7.86 3.32 ;
			RECT 5.74 2.68 7.86 3.32 ;
			RECT 6.3 2.68 6.94 9.86 ;
			RECT 6.4 2.68 6.94 11.22 ;
			RECT 6.4 10.56 7.52 11.22 ;
			RECT 7.76 4.04 8.44 9.14 ;
			RECT 7.66 8.5 9.3 9.14 ;
			RECT 10.5 1.98 11.16 3.24 ;
			RECT 9.68 2.76 11.16 3.24 ;
			RECT 9.68 2.76 10.32 5.66 ;
			RECT 9.84 2.76 10.32 11.22 ;
			RECT 9.68 10.5 10.32 11.22 ;
			RECT 12.68 3.76 14.5 4.4 ;
			RECT 12.68 3.76 13.16 8.26 ;
			RECT 11.84 7.62 13.16 8.26 ;
			RECT 11.68 1.98 12.6 2.62 ;
			RECT 11.68 1.98 12.16 4.4 ;
			RECT 10.84 3.76 12.16 4.4 ;
			RECT 10.84 3.76 11.32 9.62 ;
			RECT 10.84 8.98 14.84 9.62 ;
			RECT 13.72 8.98 14.36 11.22 ;
			RECT 16 1.98 16.86 2.62 ;
			RECT 16.38 1.98 16.86 4.62 ;
			RECT 18.74 3.36 19.38 4.62 ;
			RECT 16.38 4.14 19.38 4.62 ;
			RECT 17.44 7.42 18.12 9.06 ;
			RECT 17.44 4.14 17.92 10.04 ;
			RECT 15.6 9.56 17.92 10.04 ;
			RECT 15.6 9.56 16.08 11.22 ;
			RECT 15.16 10.5 16.08 11.22 ;
			RECT 17.38 1.98 18.38 2.8 ;
			RECT 17.38 2.32 20.38 2.8 ;
			RECT 17.38 1.98 18.02 3.62 ;
			RECT 19.9 2.32 20.38 6.5 ;
			RECT 19.34 6.02 20.38 6.5 ;
			RECT 19.34 6.02 19.82 10.06 ;
			RECT 18.92 9.42 20.56 10.06 ;
			RECT 18.44 9.58 18.92 11.22 ;
			RECT 18 10.56 18.92 11.22 ;
			RECT 21.08 1.98 22.68 2.62 ;
			RECT 21.08 1.98 21.6 6.82 ;
			RECT 21.08 5.18 23.34 6.82 ;
			RECT 20.34 7.02 21.56 8.68 ;
			RECT 21.08 1.98 21.56 11.22 ;
			RECT 19.44 10.58 21.56 11.22 ;

	END

END DFSQ

MACRO DFSHSL
	CLASS CORE ;
	FOREIGN DFSHSL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 28.8 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN C
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER MTL1 ;
			RECT 14.68 3.14 15.44 8.72 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.821 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 4.94 1.72 6.94 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.691 LAYER MTL1  ;
	END D
	PIN SB
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 9 4.92 9.68 8.94 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.851 LAYER MTL1  ;
	END SB
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 25.84 7.6 28.4 8.26 ;
			RECT 27.76 2.2 28.4 8.26 ;
			RECT 25.84 7.6 26.48 11.04 ;

		END 

		ANTENNADIFFAREA 4.598 LAYER MTL1  ;
	END Q
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 28.8 13.68 ;
			RECT 27.24 8.88 27.88 13.68 ;
			RECT 24.44 8.24 25.08 13.68 ;
			RECT 21.16 10.7 21.8 13.68 ;
			RECT 15.56 10.24 16.2 13.68 ;
			RECT 9.92 10.62 10.56 13.68 ;
			RECT 7.08 10.7 7.72 13.68 ;
			RECT 1.64 10.7 2.28 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 28.8 1.46 ;
			RECT 25.36 -0.48 26 2.84 ;
			RECT 20.08 -0.48 20.72 2.78 ;
			RECT 14.2 -0.48 14.84 2.5 ;
			RECT 9.94 -0.48 10.58 2.5 ;
			RECT 5.72 -0.48 6.36 1.78 ;
			RECT 0.42 -0.48 1.06 2.82 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 3.52 3.3 4.24 9.18 ;
			RECT 5.38 4.14 6.04 9.18 ;
			RECT 5.38 7.54 6.6 9.18 ;
			RECT 3.08 1.98 3.74 2.78 ;
			RECT 3.08 2.3 6.88 2.78 ;
			RECT 6.24 2.3 6.88 3.62 ;
			RECT 6.64 3.14 7.14 5.78 ;
			RECT 6.64 5.3 7.96 5.78 ;
			RECT 7.32 5.3 7.96 10.18 ;
			RECT 4.08 9.7 7.96 10.18 ;
			RECT 4.08 9.7 4.72 11.22 ;
			RECT 7.4 1.98 8.48 2.62 ;
			RECT 7.66 3.74 11.12 4.22 ;
			RECT 7.66 1.98 8.48 4.78 ;
			RECT 10.32 3.74 11.12 8.06 ;
			RECT 10.32 3.74 10.8 10.1 ;
			RECT 8.48 9.62 10.8 10.1 ;
			RECT 8.48 9.62 9.16 11.1 ;
			RECT 11.36 2.02 12.12 2.66 ;
			RECT 11.64 2.02 12.12 9.06 ;
			RECT 11.32 8.58 11.98 11.22 ;
			RECT 12.72 1.98 13.4 6.14 ;
			RECT 12.72 4.44 14 6.14 ;
			RECT 12.72 1.98 13.36 11.22 ;
			RECT 15.6 1.98 16.72 2.62 ;
			RECT 16 1.98 16.72 8.6 ;
			RECT 16 6.96 16.84 8.6 ;
			RECT 16 1.98 16.56 9.72 ;
			RECT 14.16 9.24 16.56 9.72 ;
			RECT 14.16 9.24 14.84 10.8 ;
			RECT 17.44 2.1 19.08 2.76 ;
			RECT 17.44 2.1 18.8 3.76 ;
			RECT 18.16 2.1 18.8 10.06 ;
			RECT 17.08 9.42 18.8 10.06 ;
			RECT 22.72 1.98 23.36 2.78 ;
			RECT 21.38 2.28 23.36 2.78 ;
			RECT 21.38 2.28 21.86 4.9 ;
			RECT 20.72 4.26 21.86 4.9 ;
			RECT 21.08 6.94 21.72 8.58 ;
			RECT 21.08 7.94 23.44 8.58 ;
			RECT 22.8 7.94 23.44 11.14 ;
			RECT 22.72 3.46 24 4.1 ;
			RECT 23.36 3.46 24 6.34 ;
			RECT 19.36 5.7 27.12 6.34 ;
			RECT 26.48 4.84 27.12 6.5 ;
			RECT 19.36 5.7 20.16 7.5 ;
			RECT 19.36 5.7 19.84 11.22 ;
			RECT 18.52 10.58 19.84 11.22 ;

	END

END DFSHSL

MACRO DFSHRL
	CLASS CORE ;
	FOREIGN DFSHRL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 33.12 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN C
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER MTL1 ;
			RECT 14.64 4.46 16.46 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.821 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 6.28 1.72 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.691 LAYER MTL1  ;
	END D
	PIN RB
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 10.24 4.18 12 4.82 ;
			RECT 10.24 4.18 11.16 9.7 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.562 LAYER MTL1  ;
	END RB
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 32.04 2.1 32.74 11.14 ;
			RECT 29.38 3.82 32.74 4.46 ;

		END 

		ANTENNADIFFAREA 6.368 LAYER MTL1  ;
	END Q
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 33.12 13.68 ;
			RECT 27.9 8.4 28.54 13.68 ;
			RECT 25.44 10.9 26.08 13.68 ;
			RECT 18.32 10.42 18.96 13.68 ;
			RECT 14.72 9.56 15.36 13.68 ;
			RECT 9.24 11.22 9.88 13.68 ;
			RECT 5.4 10.32 6.04 13.68 ;
			RECT 0.56 10.32 1.2 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 33.12 1.46 ;
			RECT 29.64 -0.48 31.28 2.7 ;
			RECT 26.08 -0.48 26.78 1.6 ;
			RECT 23.4 -0.48 24.04 2.34 ;
			RECT 17 -0.48 17.64 2.94 ;
			RECT 12.52 -0.48 13.16 2.52 ;
			RECT 9.12 -0.48 9.76 2.5 ;
			RECT 5.6 -0.48 6.24 1.78 ;
			RECT 0.4 -0.48 1.04 4.1 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 3.96 3.7 4.6 5.34 ;
			RECT 2.44 4.86 4.6 5.34 ;
			RECT 2.44 4.86 3.1 8.7 ;
			RECT 2.96 1.98 3.6 2.62 ;
			RECT 3.08 2.54 6.96 3.02 ;
			RECT 5.64 2.54 6.96 3.34 ;
			RECT 5.64 2.54 6.12 9.74 ;
			RECT 5.64 8.1 6.52 9.74 ;
			RECT 2.96 9.26 6.52 9.74 ;
			RECT 2.96 9.26 3.6 10.84 ;
			RECT 7.48 1.98 8.28 4.8 ;
			RECT 6.64 4.16 8.28 4.8 ;
			RECT 7.22 4.16 7.88 11.2 ;
			RECT 6.84 10.56 7.88 11.2 ;
			RECT 10.88 1.98 11.52 3.66 ;
			RECT 9 3.02 11.52 3.66 ;
			RECT 9 3.02 9.64 10.7 ;
			RECT 8.68 8.14 9.64 10.7 ;
			RECT 8.68 10.22 11.4 10.7 ;
			RECT 10.76 10.22 11.4 11.22 ;
			RECT 14.12 1.98 14.76 3.84 ;
			RECT 12.88 3.36 14.76 3.84 ;
			RECT 12.88 3.36 13.52 9.26 ;
			RECT 13.28 8.78 13.92 10.02 ;
			RECT 15.84 1.98 16.48 3.94 ;
			RECT 15.84 3.46 17.46 3.94 ;
			RECT 16.98 3.46 17.46 10.2 ;
			RECT 16.08 9.56 17.46 10.2 ;
			RECT 18.24 4.46 18.88 7.86 ;
			RECT 18.4 2.3 19.04 3.94 ;
			RECT 18.4 3.46 19.88 3.94 ;
			RECT 19.4 3.46 19.88 9.26 ;
			RECT 19.24 8.62 19.88 9.26 ;
			RECT 21.4 2.04 22.38 2.7 ;
			RECT 21.4 2.04 22.04 5.1 ;
			RECT 21.4 2.04 21.88 9.82 ;
			RECT 21.4 8.18 23.02 9.82 ;
			RECT 24.78 7.06 25.48 10.3 ;
			RECT 27.72 1.98 28.36 3.34 ;
			RECT 24.08 2.86 28.36 3.34 ;
			RECT 24.08 2.86 24.72 5.38 ;
			RECT 20.12 2.3 20.88 2.94 ;
			RECT 26.08 3.88 26.72 6.54 ;
			RECT 23.54 5.9 31.4 6.54 ;
			RECT 20.4 2.3 20.88 11.18 ;
			RECT 23.54 5.9 24.1 11.18 ;
			RECT 20.4 10.34 24.1 11.18 ;

	END

END DFSHRL

MACRO DFSH
	CLASS CORE ;
	FOREIGN DFSH 0 0  ;
	ORIGIN 0 0 ;
	SIZE 25.92 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN C
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER MTL1 ;
			RECT 10.12 8.56 11.78 9.2 ;
			RECT 10.48 4.96 11.12 9.2 ;
			RECT 9.76 4.96 11.12 5.6 ;
			RECT 9.76 3.58 10.4 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.821 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 0.42 6.18 1.72 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.691 LAYER MTL1  ;
	END D
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 24.5 8.58 25.52 11.22 ;
			RECT 24.88 2.16 25.52 11.22 ;
			RECT 24.8 2.16 25.52 2.8 ;

		END 

		ANTENNADIFFAREA 3.828 LAYER MTL1  ;
	END Q
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 25.92 13.68 ;
			RECT 23.04 8.58 23.68 13.68 ;
			RECT 21.16 10.7 21.8 13.68 ;
			RECT 14.24 8.58 14.88 13.68 ;
			RECT 11.28 9.92 11.92 13.68 ;
			RECT 5.32 10.7 5.96 13.68 ;
			RECT 0.44 10.7 1.08 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 25.92 1.46 ;
			RECT 23.4 -0.48 24.04 2.76 ;
			RECT 19.08 -0.48 19.72 3.7 ;
			RECT 14.28 -0.48 14.92 3.44 ;
			RECT 10.76 -0.48 11.4 2.06 ;
			RECT 5.6 -0.48 6.24 2.86 ;
			RECT 0.4 -0.48 1.04 4.42 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 3.58 4.58 4.22 9.18 ;
			RECT 2.36 8.54 4.22 9.18 ;
			RECT 2.96 2.26 3.6 2.9 ;
			RECT 3.08 2.26 3.6 3.86 ;
			RECT 3.08 3.38 6.72 3.86 ;
			RECT 5.76 3.38 6.72 4.02 ;
			RECT 5.76 3.38 6.4 9.62 ;
			RECT 5.76 3.38 6.24 10.18 ;
			RECT 2.86 9.7 6.24 10.18 ;
			RECT 2.86 9.7 3.5 11.22 ;
			RECT 7.24 2.58 8.24 3.22 ;
			RECT 7.4 2.58 8.24 5.22 ;
			RECT 7.4 2.58 8.04 11.22 ;
			RECT 6.76 10.58 8.04 11.22 ;
			RECT 9.24 1.98 9.88 3.06 ;
			RECT 8.76 2.58 11.44 3.06 ;
			RECT 10.96 2.58 11.44 3.78 ;
			RECT 10.96 3.14 12.76 3.78 ;
			RECT 8.76 2.58 9.24 10.56 ;
			RECT 8.76 6.98 9.4 10.56 ;
			RECT 8.76 9.92 10.52 10.56 ;
			RECT 12.52 1.98 13.76 2.62 ;
			RECT 13.28 1.98 13.76 6.22 ;
			RECT 12.72 5.58 14.38 6.22 ;
			RECT 12.72 5.58 13.36 10.12 ;
			RECT 15.68 2.8 16.32 11.22 ;
			RECT 20.52 8.54 22.16 9.18 ;
			RECT 20.52 8.54 21.16 10.18 ;
			RECT 20.52 1.98 22.36 2.62 ;
			RECT 20.52 1.98 21.16 6.58 ;
			RECT 21.72 3.44 24.36 4.08 ;
			RECT 21.72 3.44 22.2 8.02 ;
			RECT 17.08 7.38 24.2 8.02 ;
			RECT 17.08 2.8 17.72 11.22 ;
			RECT 17.08 10.58 19.16 11.22 ;

	END

END DFSH

MACRO DFMSLQ
	CLASS CORE ;
	FOREIGN DFMSLQ 0 0  ;
	ORIGIN 0 0 ;
	SIZE 36 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN C
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER MTL1 ;
			RECT 25.44 6.28 26.08 9.04 ;
			RECT 23.44 6.28 26.08 6.92 ;
			RECT 23.44 4.96 24.84 6.92 ;
			RECT 24.08 3.54 24.84 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.821 LAYER MTL1  ;
	END C
	PIN D0
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.42 2.48 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.662 LAYER MTL1  ;
	END D0
	PIN D1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 6.6 7.6 8.24 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.662 LAYER MTL1  ;
	END D1
	PIN S1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.31 LAYER MTL1  ;
	END S1
	PIN SB
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 16 9.22 17.64 9.86 ;
			RECT 16.24 3.14 16.96 4.78 ;
			RECT 16.24 3.14 16.88 9.86 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.57 LAYER MTL1  ;
	END SB
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 34.96 1.98 35.6 11.22 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END Q
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 36 13.68 ;
			RECT 33.56 9.12 34.2 13.68 ;
			RECT 32.12 10.58 32.76 13.68 ;
			RECT 26.32 10.68 26.96 13.68 ;
			RECT 21.08 10.32 21.72 13.68 ;
			RECT 18 10.58 18.64 13.68 ;
			RECT 15.36 10.58 16 13.68 ;
			RECT 12.56 10.7 13.2 13.68 ;
			RECT 6.64 10.7 7.28 13.68 ;
			RECT 1.8 10.58 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 36 1.46 ;
			RECT 33.56 -0.48 34.2 2.66 ;
			RECT 28.02 -0.48 28.66 1.8 ;
			RECT 23.2 -0.48 23.84 2.54 ;
			RECT 16.96 -0.48 17.6 2.62 ;
			RECT 12.88 -0.48 13.52 2.62 ;
			RECT 6.88 -0.48 7.52 2.26 ;
			RECT 1 -0.48 1.64 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1 3.14 4.24 3.9 ;
			RECT 3.6 3.14 4.24 4.78 ;
			RECT 3.6 4.3 5.42 4.78 ;
			RECT 4.76 4.3 5.42 9.18 ;
			RECT 3 8.7 5.42 9.18 ;
			RECT 3 8.7 3.48 10.06 ;
			RECT 0.4 9.58 3.48 10.06 ;
			RECT 0.4 9.58 1.04 11.22 ;
			RECT 4.24 9.7 9.24 10.18 ;
			RECT 4.24 9.7 4.88 11.22 ;
			RECT 8.6 9.7 9.24 11.22 ;
			RECT 4.24 1.98 5.52 2.62 ;
			RECT 5 1.98 5.52 3.26 ;
			RECT 8.6 1.98 9.24 3.26 ;
			RECT 5 2.78 9.24 3.26 ;
			RECT 9.76 3.14 11.24 4.78 ;
			RECT 9.76 3.14 10.24 9.18 ;
			RECT 9.48 7.54 10.24 9.18 ;
			RECT 10.24 1.98 12.3 2.62 ;
			RECT 11.8 1.98 12.3 3.8 ;
			RECT 11.8 3.14 13.88 3.8 ;
			RECT 11.8 9.22 13.56 9.86 ;
			RECT 11.8 1.98 12.28 10.18 ;
			RECT 10 9.7 12.28 10.18 ;
			RECT 10 9.7 10.64 11.22 ;
			RECT 14.32 1.98 14.96 2.62 ;
			RECT 14.4 1.98 14.88 5 ;
			RECT 12.8 4.52 14.56 5.16 ;
			RECT 14.08 4.52 14.56 11.22 ;
			RECT 13.06 7.84 14.7 8.48 ;
			RECT 14.08 7.84 14.7 11.22 ;
			RECT 13.96 10.58 14.7 11.22 ;
			RECT 18.12 1.98 20 2.62 ;
			RECT 18.12 1.98 18.6 6.18 ;
			RECT 18.12 5.54 20.08 6.18 ;
			RECT 19.16 5.54 19.64 10.7 ;
			RECT 19.16 10.06 20.28 10.7 ;
			RECT 21.6 3.54 23.34 4.18 ;
			RECT 21.6 3.54 22.08 8.54 ;
			RECT 21.6 7.9 22.24 8.54 ;
			RECT 20.6 1.98 21.44 2.62 ;
			RECT 19.12 3.14 21.08 4.78 ;
			RECT 23.48 8.26 24.6 8.9 ;
			RECT 20.6 1.98 21.08 9.54 ;
			RECT 20.16 8.9 21.08 9.54 ;
			RECT 20.16 9.06 24.12 9.54 ;
			RECT 23.48 8.26 24.12 11.22 ;
			RECT 24.72 1.98 25.86 2.62 ;
			RECT 25.38 1.98 25.86 3.96 ;
			RECT 25.38 3.32 27.08 3.96 ;
			RECT 26.6 8.4 27.48 9.06 ;
			RECT 26.6 3.32 27.08 10.04 ;
			RECT 24.92 9.56 27.08 10.04 ;
			RECT 24.92 9.56 25.6 11.22 ;
			RECT 26.38 1.98 27.02 2.8 ;
			RECT 26.38 2.32 29.02 2.8 ;
			RECT 27.68 4.54 29.02 5.18 ;
			RECT 28.54 2.32 29.02 10.06 ;
			RECT 28.54 9.42 30.44 10.06 ;
			RECT 28.16 9.58 28.64 11.22 ;
			RECT 27.72 10.58 28.64 11.22 ;
			RECT 30.68 1.98 31.56 2.62 ;
			RECT 29.54 6.9 31.56 8.54 ;
			RECT 31.04 1.98 31.56 11.22 ;
			RECT 29.16 10.58 31.56 11.22 ;
			RECT 32.12 3.66 33.36 4.3 ;
			RECT 32.12 5.18 32.84 6.82 ;
			RECT 32.12 3.66 32.76 9.74 ;

	END

END DFMSLQ

MACRO DFMRLSLQ
	CLASS CORE ;
	FOREIGN DFMRLSLQ 0 0  ;
	ORIGIN 0 0 ;
	SIZE 41.76 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN C
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER MTL1 ;
			RECT 31.16 6.28 31.8 9.04 ;
			RECT 29.2 7.6 31.8 8.24 ;
			RECT 29.62 6.28 31.8 8.24 ;
			RECT 29.62 3.76 30.26 8.24 ;
			RECT 29.2 6.28 31.8 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.821 LAYER MTL1  ;
	END C
	PIN D0
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.42 2.48 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.691 LAYER MTL1  ;
	END D0
	PIN D1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 6.6 7.6 8.24 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.691 LAYER MTL1  ;
	END D1
	PIN S1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.339 LAYER MTL1  ;
	END S1
	PIN RB
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 19.28 4.54 19.96 5.18 ;
			RECT 18.34 6.28 19.76 8.24 ;
			RECT 19.28 4.54 19.76 8.24 ;
			RECT 18.34 6.28 19.16 9.56 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.562 LAYER MTL1  ;
	END RB
	PIN SB
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 21.52 8.9 23.2 9.54 ;
			RECT 22.72 5.54 23.2 9.54 ;
			RECT 21.48 5.54 23.2 6.18 ;
			RECT 11.8 3.14 13.88 3.8 ;
			RECT 11.8 9.46 13.56 10.14 ;
			RECT 11.8 7.6 12.56 10.14 ;
			RECT 11.8 6.28 12.56 6.92 ;
			RECT 11.8 3.14 12.28 10.14 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.872 LAYER MTL1  ;
	END SB
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 40.72 1.98 41.36 11.22 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END Q
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 41.76 13.68 ;
			RECT 39.32 9.26 39.96 13.68 ;
			RECT 37.88 10.58 38.52 13.68 ;
			RECT 32.08 10.68 32.72 13.68 ;
			RECT 26.8 10.32 27.44 13.68 ;
			RECT 22.44 11.06 23.08 13.68 ;
			RECT 17.52 10.58 18.16 13.68 ;
			RECT 12.56 11.66 13.2 13.68 ;
			RECT 6.64 10.7 7.28 13.68 ;
			RECT 1.8 10.58 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 41.76 1.46 ;
			RECT 39.32 -0.48 39.96 2.66 ;
			RECT 33.78 -0.48 34.42 1.8 ;
			RECT 28.76 -0.48 29.4 2.54 ;
			RECT 20.6 -0.48 21.24 2.5 ;
			RECT 12.88 -0.48 13.52 2.58 ;
			RECT 6.88 -0.48 7.52 2.26 ;
			RECT 1 -0.48 1.64 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1 3.14 4.24 3.9 ;
			RECT 3.6 3.14 4.24 4.78 ;
			RECT 3.6 4.14 5.4 4.78 ;
			RECT 4.76 4.14 5.4 9.04 ;
			RECT 3 8.56 5.4 9.04 ;
			RECT 3 8.56 3.48 10.06 ;
			RECT 0.4 9.58 3.48 10.06 ;
			RECT 0.4 9.58 1.04 11.22 ;
			RECT 4.24 9.7 8.36 10.18 ;
			RECT 7.88 9.7 8.36 11.22 ;
			RECT 4.24 9.7 4.88 11.22 ;
			RECT 7.88 10.58 9.24 11.22 ;
			RECT 4.24 1.98 5.52 2.62 ;
			RECT 5 1.98 5.52 3.26 ;
			RECT 8.6 1.98 9.24 3.26 ;
			RECT 5 2.78 9.24 3.26 ;
			RECT 9.64 3.98 10.28 9.44 ;
			RECT 9.56 7.78 10.28 9.44 ;
			RECT 15.8 2.98 16.44 5 ;
			RECT 12.8 4.52 16.44 5 ;
			RECT 12.8 4.52 14.76 5.16 ;
			RECT 14.28 4.52 14.76 8.54 ;
			RECT 14.48 7.9 15.12 10.14 ;
			RECT 10.24 1.98 11.28 2.62 ;
			RECT 16.96 3.14 17.6 3.78 ;
			RECT 16.96 3.14 17.44 9.7 ;
			RECT 15.64 9.06 17.44 9.7 ;
			RECT 10.8 1.98 11.28 11.14 ;
			RECT 10 10.58 11.28 11.14 ;
			RECT 15.64 9.06 16.12 11.14 ;
			RECT 10 10.66 16.12 11.14 ;
			RECT 10 10.58 10.64 11.22 ;
			RECT 14.28 1.98 17.96 2.46 ;
			RECT 14.28 1.98 14.92 2.62 ;
			RECT 17.32 1.98 17.96 2.62 ;
			RECT 18.96 1.98 19.6 4.02 ;
			RECT 18.12 3.54 23 4.02 ;
			RECT 22.52 3.54 23 4.78 ;
			RECT 22.52 4.14 23.16 4.78 ;
			RECT 18.12 3.54 18.6 5.18 ;
			RECT 17.96 4.54 18.6 5.18 ;
			RECT 20.48 3.54 20.96 9.54 ;
			RECT 19.68 8.9 20.96 9.54 ;
			RECT 19.68 8.9 20.2 11.22 ;
			RECT 19.08 10.58 20.2 11.22 ;
			RECT 23.52 2.98 24.2 3.62 ;
			RECT 23.72 5.54 25.36 6.18 ;
			RECT 23.72 2.98 24.2 10.54 ;
			RECT 20.92 10.06 25.48 10.54 ;
			RECT 20.92 10.06 21.56 11.22 ;
			RECT 24.84 10.06 25.48 11.22 ;
			RECT 22 1.98 25.56 2.46 ;
			RECT 22 1.98 22.64 2.62 ;
			RECT 24.92 1.98 25.56 3.34 ;
			RECT 27.2 3.76 28.9 4.4 ;
			RECT 27.2 3.76 27.68 8.54 ;
			RECT 27.2 7.9 27.84 8.54 ;
			RECT 26.2 1.98 27 2.62 ;
			RECT 24.72 3.98 26.68 4.62 ;
			RECT 26.2 1.98 26.68 9.54 ;
			RECT 25.84 8.9 26.68 9.54 ;
			RECT 29.24 8.9 30.36 9.54 ;
			RECT 25.84 9.06 30.36 9.54 ;
			RECT 29.2 9.06 29.84 11.22 ;
			RECT 30.4 1.98 31.26 2.62 ;
			RECT 30.78 1.98 31.26 4.62 ;
			RECT 33.14 3.36 33.78 4.62 ;
			RECT 30.78 4.14 33.78 4.62 ;
			RECT 32.8 7.4 33.6 9.06 ;
			RECT 32.8 4.14 33.28 10.04 ;
			RECT 30.88 9.56 33.28 10.04 ;
			RECT 30.88 9.56 31.36 11.22 ;
			RECT 30.64 10.5 31.36 11.22 ;
			RECT 31.78 1.98 32.78 2.8 ;
			RECT 31.78 2.32 34.78 2.8 ;
			RECT 31.78 1.98 32.42 3.62 ;
			RECT 34.3 2.32 34.78 10.06 ;
			RECT 34.3 9.42 36.2 10.06 ;
			RECT 33.92 9.58 34.4 11.22 ;
			RECT 33.48 10.58 34.4 11.22 ;
			RECT 35.3 1.98 37.08 2.62 ;
			RECT 35.3 1.98 35.94 8.9 ;
			RECT 35.3 8.42 37.2 8.9 ;
			RECT 36.72 8.42 37.2 11.22 ;
			RECT 34.92 10.58 37.2 11.22 ;
			RECT 36.46 3.66 39.12 4.3 ;
			RECT 36.46 3.66 36.94 7.5 ;
			RECT 36.46 7.02 38.56 7.5 ;
			RECT 37.84 7.02 38.56 9.74 ;

	END

END DFMRLSLQ

MACRO DFMRLQ
	CLASS CORE ;
	FOREIGN DFMRLQ 0 0  ;
	ORIGIN 0 0 ;
	SIZE 38.88 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN C
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER MTL1 ;
			RECT 28.28 6.28 28.92 9.04 ;
			RECT 26.32 7.6 28.92 8.24 ;
			RECT 26.74 6.28 28.92 8.24 ;
			RECT 26.74 3.76 27.38 8.24 ;
			RECT 26.32 6.28 28.92 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.821 LAYER MTL1  ;
	END C
	PIN D0
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.42 2.48 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.691 LAYER MTL1  ;
	END D0
	PIN D1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 6.6 7.6 8.24 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.691 LAYER MTL1  ;
	END D1
	PIN S1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.339 LAYER MTL1  ;
	END S1
	PIN RB
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 17.56 8.9 19.76 9.56 ;
			RECT 19.12 3.14 19.76 9.56 ;
			RECT 18.6 3.14 19.76 4.78 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.562 LAYER MTL1  ;
	END RB
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 37.84 1.98 38.48 11.22 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END Q
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 38.88 13.68 ;
			RECT 36.44 9.1 37.08 13.68 ;
			RECT 35 10.58 35.64 13.68 ;
			RECT 29.2 10.68 29.84 13.68 ;
			RECT 23.92 10.74 24.56 13.68 ;
			RECT 19.56 10.38 20.2 13.68 ;
			RECT 15.88 11.22 16.52 13.68 ;
			RECT 12.04 10.7 12.68 13.68 ;
			RECT 6.64 10.7 7.28 13.68 ;
			RECT 1.8 10.58 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 38.88 1.46 ;
			RECT 36.44 -0.48 37.08 2.66 ;
			RECT 30.9 -0.48 31.54 1.8 ;
			RECT 25.88 -0.48 26.52 2.82 ;
			RECT 22.02 -0.48 22.68 2.62 ;
			RECT 19.24 -0.48 19.88 2.62 ;
			RECT 16.16 -0.48 16.8 2.14 ;
			RECT 12.88 -0.48 13.52 1.78 ;
			RECT 6.88 -0.48 7.52 2.26 ;
			RECT 1 -0.48 1.64 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1 3.14 4.24 3.9 ;
			RECT 3.6 3.14 4.24 4.78 ;
			RECT 3.6 4.3 5.4 4.78 ;
			RECT 4.76 4.3 5.4 9.14 ;
			RECT 3 8.64 5.4 9.14 ;
			RECT 3 8.64 3.48 10.06 ;
			RECT 0.4 9.58 3.48 10.06 ;
			RECT 0.4 9.58 1.04 11.22 ;
			RECT 4.24 9.7 8.84 10.18 ;
			RECT 4.24 9.7 4.88 11.22 ;
			RECT 8.2 9.7 8.84 11.22 ;
			RECT 4.24 1.98 5.52 2.62 ;
			RECT 5 1.98 5.52 3.26 ;
			RECT 8.58 1.98 9.22 3.26 ;
			RECT 5 2.78 9.22 3.26 ;
			RECT 10.84 3.3 11.48 9.18 ;
			RECT 9.08 7.54 11.48 9.18 ;
			RECT 14.52 1.98 15.16 2.78 ;
			RECT 13.16 2.3 15.16 2.78 ;
			RECT 13.16 2.3 13.8 8.34 ;
			RECT 15.32 7.7 15.96 10.7 ;
			RECT 13.48 10.22 15.96 10.7 ;
			RECT 13.48 10.22 14.18 10.86 ;
			RECT 10.22 1.98 10.9 2.78 ;
			RECT 10.22 2.3 12.48 2.78 ;
			RECT 15.68 2.66 16.32 3.78 ;
			RECT 14.32 3.3 16.32 3.78 ;
			RECT 12 9.06 14.8 9.7 ;
			RECT 14.32 3.3 14.8 9.7 ;
			RECT 12 2.3 12.48 10.18 ;
			RECT 9.6 9.7 12.48 10.18 ;
			RECT 9.6 9.7 10.24 11.22 ;
			RECT 17.32 1.98 18.24 2.62 ;
			RECT 17.32 1.98 17.8 4.94 ;
			RECT 15.48 4.3 17.8 4.94 ;
			RECT 16.48 4.3 16.96 10.7 ;
			RECT 16.48 10.22 19.04 10.7 ;
			RECT 17.4 10.22 19.04 11.22 ;
			RECT 20.64 1.98 21.5 2.62 ;
			RECT 21.02 1.98 21.5 3.62 ;
			RECT 21.02 3.14 22.28 3.62 ;
			RECT 21.64 3.14 22.28 5.4 ;
			RECT 21.76 3.14 22.28 10.92 ;
			RECT 21.76 10.26 22.6 10.92 ;
			RECT 24.2 3.76 26.02 4.4 ;
			RECT 24.2 3.76 24.68 8.38 ;
			RECT 24.16 7.7 24.8 8.38 ;
			RECT 23.2 1.98 24.12 2.62 ;
			RECT 23.2 1.98 23.68 4.38 ;
			RECT 22.92 3.74 23.4 9.74 ;
			RECT 26.36 8.9 27.48 9.54 ;
			RECT 22.92 9.08 26.96 9.74 ;
			RECT 26.32 9.08 26.96 11.22 ;
			RECT 27.52 1.98 28.38 2.62 ;
			RECT 27.9 1.98 28.38 4.62 ;
			RECT 30.26 3.36 30.9 4.62 ;
			RECT 27.9 4.14 30.9 4.62 ;
			RECT 29.92 7.42 30.72 9.06 ;
			RECT 29.92 4.14 30.4 10.04 ;
			RECT 28 9.56 30.4 10.04 ;
			RECT 28 9.56 28.48 11.22 ;
			RECT 27.76 10.5 28.48 11.22 ;
			RECT 28.9 1.98 29.9 2.8 ;
			RECT 28.9 2.32 31.9 2.8 ;
			RECT 28.9 1.98 29.54 3.62 ;
			RECT 31.42 2.32 31.9 10.06 ;
			RECT 31.42 8.9 32.12 10.06 ;
			RECT 31.04 9.58 31.52 11.22 ;
			RECT 30.6 10.58 31.52 11.22 ;
			RECT 32.64 1.98 34.2 2.62 ;
			RECT 32.42 6.22 33.12 7.86 ;
			RECT 32.64 1.98 33.12 11.22 ;
			RECT 32.04 10.58 33.12 11.22 ;
			RECT 33.64 3.66 36.24 4.3 ;
			RECT 33.64 3.66 34.12 7.52 ;
			RECT 33.64 7.02 35.68 7.52 ;
			RECT 34.96 7.02 35.68 9.74 ;

	END

END DFMRLQ

MACRO DFMQ
	CLASS CORE ;
	FOREIGN DFMQ 0 0  ;
	ORIGIN 0 0 ;
	SIZE 33.12 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN C
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER MTL1 ;
			RECT 22 7.6 24.08 8.24 ;
			RECT 22.42 6.28 24.08 8.24 ;
			RECT 23.24 6.28 23.88 9.04 ;
			RECT 22.42 3.76 23.06 8.24 ;
			RECT 22 6.28 24.08 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.821 LAYER MTL1  ;
	END C
	PIN D0
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.42 2.48 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.634 LAYER MTL1  ;
	END D0
	PIN D1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 6.6 7.6 8.24 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.634 LAYER MTL1  ;
	END D1
	PIN S1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.282 LAYER MTL1  ;
	END S1
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 32.08 1.98 32.72 11.22 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END Q
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 33.12 13.68 ;
			RECT 29.28 10.58 31.32 13.68 ;
			RECT 30.68 9.1 31.32 13.68 ;
			RECT 23.8 10.68 24.44 13.68 ;
			RECT 18.52 10.14 19.16 13.68 ;
			RECT 15.48 10.38 16.12 13.68 ;
			RECT 12.44 10.7 13.08 13.68 ;
			RECT 6.6 10.7 7.24 13.68 ;
			RECT 1.8 10.58 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 33.12 1.46 ;
			RECT 30.68 -0.48 31.32 2.26 ;
			RECT 26.58 -0.48 27.22 1.8 ;
			RECT 21.56 -0.48 22.2 2.82 ;
			RECT 16.06 -0.48 16.7 2.14 ;
			RECT 12.98 -0.48 13.62 1.78 ;
			RECT 6.88 -0.48 7.52 2.26 ;
			RECT 1 -0.48 1.64 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1 3.14 4.24 3.9 ;
			RECT 3 3.14 4.24 4.78 ;
			RECT 3 7.54 5.38 9.18 ;
			RECT 3 3.14 3.48 10.06 ;
			RECT 0.4 9.58 3.48 10.06 ;
			RECT 0.4 9.58 1.04 11.22 ;
			RECT 4.2 9.7 9.24 10.18 ;
			RECT 4.2 9.7 4.84 11.22 ;
			RECT 8.6 9.7 9.24 11.22 ;
			RECT 4.24 1.98 5.52 2.62 ;
			RECT 5 1.98 5.52 3.26 ;
			RECT 8.6 1.98 9.24 3.26 ;
			RECT 5 2.78 9.24 3.26 ;
			RECT 10.68 3.3 11.32 8.02 ;
			RECT 9.48 7.54 11.32 8.02 ;
			RECT 9.48 7.54 10.12 9.18 ;
			RECT 10.32 1.98 11 2.78 ;
			RECT 10.32 2.3 12.42 2.78 ;
			RECT 11.94 4.04 12.98 5.68 ;
			RECT 11.94 2.3 12.42 10.18 ;
			RECT 10 9.7 12.42 10.18 ;
			RECT 10 9.7 10.64 11.22 ;
			RECT 14.42 1.98 15.06 3.32 ;
			RECT 12.94 2.68 15.06 3.32 ;
			RECT 13.5 2.68 14.14 9.7 ;
			RECT 13.6 2.68 14.14 11.22 ;
			RECT 13.6 10.56 14.72 11.22 ;
			RECT 14.96 4.04 15.64 9.7 ;
			RECT 17.7 1.98 18.36 3.24 ;
			RECT 16.88 2.76 18.36 3.24 ;
			RECT 16.88 2.76 17.52 11.22 ;
			RECT 19.88 3.76 21.7 4.4 ;
			RECT 19.88 3.76 20.36 8.26 ;
			RECT 19.04 7.62 20.36 8.26 ;
			RECT 18.88 1.98 19.8 2.62 ;
			RECT 18.88 1.98 19.36 4.4 ;
			RECT 18.04 3.76 19.36 4.4 ;
			RECT 18.04 3.76 18.52 9.62 ;
			RECT 18.04 8.98 22.04 9.62 ;
			RECT 20.92 8.98 21.56 11.22 ;
			RECT 23.2 1.98 24.06 2.62 ;
			RECT 23.58 1.98 24.06 4.62 ;
			RECT 25.94 3.36 26.58 4.62 ;
			RECT 23.58 4.14 26.58 4.62 ;
			RECT 24.64 7.42 25.32 9.06 ;
			RECT 24.64 4.14 25.12 10.04 ;
			RECT 22.8 9.56 25.12 10.04 ;
			RECT 22.8 9.56 23.28 11.22 ;
			RECT 22.36 10.5 23.28 11.22 ;
			RECT 24.58 1.98 25.58 2.8 ;
			RECT 24.58 2.32 27.58 2.8 ;
			RECT 24.58 1.98 25.22 3.62 ;
			RECT 27.1 2.32 27.58 5.62 ;
			RECT 26.08 5.14 27.58 5.62 ;
			RECT 26.08 5.14 26.56 10.06 ;
			RECT 26.08 9.42 27.76 10.06 ;
			RECT 25.64 9.58 26.12 11.22 ;
			RECT 25.2 10.56 26.12 11.22 ;
			RECT 28.28 1.98 29.88 2.62 ;
			RECT 28.28 1.98 28.8 6.82 ;
			RECT 28.28 5.18 30.08 6.82 ;
			RECT 27.08 6.42 28.76 8.06 ;
			RECT 28.28 1.98 28.76 11.22 ;
			RECT 26.64 10.58 28.76 11.22 ;

	END

END DFMQ

MACRO DFMHSL
	CLASS CORE ;
	FOREIGN DFMHSL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 36 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN C
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER MTL1 ;
			RECT 21.88 3.14 22.64 8.72 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.821 LAYER MTL1  ;
	END C
	PIN D0
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.42 2.48 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.734 LAYER MTL1  ;
	END D0
	PIN D1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 6.6 7.6 8.24 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.734 LAYER MTL1  ;
	END D1
	PIN S1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.382 LAYER MTL1  ;
	END S1
	PIN SB
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 16.24 3.74 16.96 4.38 ;
			RECT 15.08 8.78 16.88 9.42 ;
			RECT 16.24 3.64 16.88 9.42 ;
			RECT 15.08 8.78 15.72 9.86 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.779 LAYER MTL1  ;
	END SB
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 33.04 7.6 35.6 8.26 ;
			RECT 34.96 2.2 35.6 8.26 ;
			RECT 33.04 7.6 33.68 11.04 ;

		END 

		ANTENNADIFFAREA 4.598 LAYER MTL1  ;
	END Q
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 36 13.68 ;
			RECT 34.44 8.88 35.08 13.68 ;
			RECT 31.64 8.24 32.28 13.68 ;
			RECT 28.36 10.7 29 13.68 ;
			RECT 22.76 10.24 23.4 13.68 ;
			RECT 15.46 10.58 16.1 13.68 ;
			RECT 12.56 10.7 13.2 13.68 ;
			RECT 6.64 10.7 7.28 13.68 ;
			RECT 1.8 10.58 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 36 1.46 ;
			RECT 32.56 -0.48 33.2 2.84 ;
			RECT 27.28 -0.48 27.92 2.78 ;
			RECT 21.4 -0.48 22.04 2.5 ;
			RECT 16.96 -0.48 17.6 2.62 ;
			RECT 12.88 -0.48 13.52 2.62 ;
			RECT 6.88 -0.48 7.52 2.26 ;
			RECT 1 -0.48 1.64 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1 3.14 4.24 3.9 ;
			RECT 3.6 3.14 4.24 4.78 ;
			RECT 3.6 4.3 5.42 4.78 ;
			RECT 4.76 4.3 5.42 9.18 ;
			RECT 3 8.7 5.42 9.18 ;
			RECT 3 8.7 3.48 10.06 ;
			RECT 0.4 9.58 3.48 10.06 ;
			RECT 0.4 9.58 1.04 11.22 ;
			RECT 4.24 9.7 9.24 10.18 ;
			RECT 4.24 9.7 4.88 11.22 ;
			RECT 8.6 9.7 9.24 11.22 ;
			RECT 4.24 1.98 5.52 2.62 ;
			RECT 5 1.98 5.52 3.26 ;
			RECT 8.6 1.98 9.24 3.26 ;
			RECT 5 2.78 9.24 3.26 ;
			RECT 9.76 3.14 11.24 4.78 ;
			RECT 9.76 3.14 10.24 9.18 ;
			RECT 9.48 7.54 10.24 9.18 ;
			RECT 10.24 1.98 12.24 2.62 ;
			RECT 11.76 3.14 13.88 3.8 ;
			RECT 11.76 9.22 13.56 9.86 ;
			RECT 11.76 1.98 12.24 10.18 ;
			RECT 10 9.7 12.24 10.18 ;
			RECT 10 9.7 10.64 11.22 ;
			RECT 14.32 1.98 14.96 2.62 ;
			RECT 14.4 1.98 14.88 5.22 ;
			RECT 12.92 4.74 14.56 5.38 ;
			RECT 12.92 7.78 14.56 8.42 ;
			RECT 14.08 4.74 14.56 11.22 ;
			RECT 13.96 10.58 14.6 11.22 ;
			RECT 18.36 1.98 19 8.06 ;
			RECT 17.4 7.44 19 8.06 ;
			RECT 17.4 7.44 18.04 11.22 ;
			RECT 19.76 1.98 20.4 9.22 ;
			RECT 18.8 8.58 20.4 9.22 ;
			RECT 18.8 8.58 19.44 11.22 ;
			RECT 22.8 1.98 23.92 2.62 ;
			RECT 23.2 1.98 23.92 8.46 ;
			RECT 23.2 6.82 24.04 8.46 ;
			RECT 23.2 1.98 23.76 9.72 ;
			RECT 21.36 9.24 23.76 9.72 ;
			RECT 21.36 9.24 22.04 10.8 ;
			RECT 24.64 2.1 26.28 2.76 ;
			RECT 24.64 2.1 26 3.76 ;
			RECT 25.36 2.1 26 10.06 ;
			RECT 24.28 9.42 26 10.06 ;
			RECT 29.92 1.98 30.56 2.78 ;
			RECT 28.58 2.28 30.56 2.78 ;
			RECT 28.58 2.28 29.06 4.9 ;
			RECT 27.92 4.26 29.06 4.9 ;
			RECT 28.28 6.94 28.92 8.58 ;
			RECT 28.28 7.94 30.64 8.58 ;
			RECT 30 7.94 30.64 11.14 ;
			RECT 29.92 3.46 31.2 4.1 ;
			RECT 30.56 3.46 31.2 6.34 ;
			RECT 26.56 5.7 34.32 6.34 ;
			RECT 33.68 4.84 34.32 6.5 ;
			RECT 26.56 5.7 27.36 7.5 ;
			RECT 26.56 5.7 27.04 11.22 ;
			RECT 25.72 10.58 27.04 11.22 ;

	END

END DFMHSL

MACRO DFMHRL
	CLASS CORE ;
	FOREIGN DFMHRL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 38.88 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN C
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER MTL1 ;
			RECT 20.4 4.46 22.22 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.821 LAYER MTL1  ;
	END C
	PIN D0
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.42 2.48 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.734 LAYER MTL1  ;
	END D0
	PIN D1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 6.6 6.88 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.734 LAYER MTL1  ;
	END D1
	PIN S1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.382 LAYER MTL1  ;
	END S1
	PIN RB
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 16.84 6.28 18.32 9.7 ;
			RECT 16.84 4.18 17.52 9.7 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.562 LAYER MTL1  ;
	END RB
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 37.8 2.1 38.5 11.14 ;
			RECT 35.34 3.82 38.5 4.46 ;

		END 

		ANTENNADIFFAREA 6.368 LAYER MTL1  ;
	END Q
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 38.88 13.68 ;
			RECT 33.66 8.4 34.3 13.68 ;
			RECT 31.2 10.9 31.84 13.68 ;
			RECT 24.08 10.42 24.72 13.68 ;
			RECT 20.48 9.56 21.12 13.68 ;
			RECT 15.84 11.22 16.48 13.68 ;
			RECT 12 10.4 12.64 13.68 ;
			RECT 6.64 10.7 7.28 13.68 ;
			RECT 1.8 10.58 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 38.88 1.46 ;
			RECT 35.4 -0.48 37.04 2.7 ;
			RECT 31.88 -0.48 32.58 1.9 ;
			RECT 29.24 -0.48 29.88 2.34 ;
			RECT 23.36 -0.48 24 2.94 ;
			RECT 19.64 -0.48 20.28 2.52 ;
			RECT 16.12 -0.48 16.76 2.62 ;
			RECT 13.32 -0.48 13.96 2.62 ;
			RECT 6.88 -0.48 7.52 2.26 ;
			RECT 1 -0.48 1.64 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1 3.14 4.24 3.9 ;
			RECT 3.6 3.14 4.24 4.78 ;
			RECT 3.6 4.3 5.4 4.78 ;
			RECT 4.76 4.3 5.4 9.14 ;
			RECT 3 8.64 5.4 9.14 ;
			RECT 3 8.64 3.48 10.06 ;
			RECT 0.4 9.58 3.48 10.06 ;
			RECT 0.4 9.58 1.04 11.22 ;
			RECT 4.24 9.7 8.72 10.18 ;
			RECT 8.08 9.7 8.72 10.92 ;
			RECT 4.24 9.7 4.88 11.22 ;
			RECT 4.24 1.98 5.52 2.62 ;
			RECT 5 1.98 5.52 3.62 ;
			RECT 5 3.14 11.8 3.62 ;
			RECT 11.16 3.14 11.8 3.78 ;
			RECT 7.52 4.14 8.16 5.8 ;
			RECT 7.52 5.22 12.12 5.8 ;
			RECT 11.48 5.22 12.12 8.42 ;
			RECT 9.52 1.98 12.8 2.62 ;
			RECT 12.32 1.98 12.8 3.78 ;
			RECT 12.32 3.14 13.48 3.78 ;
			RECT 12.82 3.14 13.48 9.78 ;
			RECT 9.48 9.14 13.48 9.78 ;
			RECT 9.48 9.14 10.12 10.58 ;
			RECT 14.48 1.98 15.36 2.62 ;
			RECT 14.48 1.98 15 3.66 ;
			RECT 14 3.14 14.64 11.2 ;
			RECT 13.44 10.56 14.64 11.2 ;
			RECT 17.56 1.98 18.2 3.66 ;
			RECT 15.52 3.14 18.2 3.66 ;
			RECT 15.52 3.14 16.16 10.7 ;
			RECT 15.52 10.22 18.04 10.7 ;
			RECT 17.4 10.22 18.04 11.22 ;
			RECT 21.04 1.98 21.68 3.84 ;
			RECT 19.16 3.36 21.68 3.84 ;
			RECT 19.16 3.36 19.8 10.02 ;
			RECT 19 9.26 19.8 10.02 ;
			RECT 22.2 1.98 22.84 3.94 ;
			RECT 22.74 3.46 23.22 10.2 ;
			RECT 21.84 9.56 23.22 10.2 ;
			RECT 24 3.76 24.64 7.86 ;
			RECT 24.76 2.3 25.64 2.94 ;
			RECT 25.16 2.3 25.64 9.26 ;
			RECT 25 8.62 25.64 9.26 ;
			RECT 27.32 2.04 28.24 2.7 ;
			RECT 27.32 2.04 27.8 5.1 ;
			RECT 27.16 3.46 27.64 9.82 ;
			RECT 27.16 8.18 28.78 9.82 ;
			RECT 30.54 7.06 31.24 10.3 ;
			RECT 33.52 1.98 34.16 3.34 ;
			RECT 29.88 2.86 34.16 3.34 ;
			RECT 29.88 2.86 30.52 5.38 ;
			RECT 26.16 2.3 26.8 2.94 ;
			RECT 31.88 3.88 32.52 6.54 ;
			RECT 29.3 5.9 37.16 6.54 ;
			RECT 26.16 2.3 26.64 11.18 ;
			RECT 29.3 5.9 29.86 11.18 ;
			RECT 26.16 10.34 29.86 11.18 ;

	END

END DFMHRL

MACRO DFMH
	CLASS CORE ;
	FOREIGN DFMH 0 0  ;
	ORIGIN 0 0 ;
	SIZE 33.12 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN C
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER MTL1 ;
			RECT 17.32 8.56 18.98 9.2 ;
			RECT 17.68 4.96 18.32 9.2 ;
			RECT 16.96 4.96 18.32 5.6 ;
			RECT 16.96 3.58 17.6 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.821 LAYER MTL1  ;
	END C
	PIN D0
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 2.84 7.2 3.92 8.86 ;
			RECT 3.28 4.42 3.92 8.86 ;
			RECT 2.22 4.42 3.92 5.06 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.691 LAYER MTL1  ;
	END D0
	PIN D1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 7.1 4.96 8.24 7.06 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.691 LAYER MTL1  ;
	END D1
	PIN S1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 4.96 1.5 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.339 LAYER MTL1  ;
	END S1
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 31.7 8.58 32.72 11.22 ;
			RECT 32.08 2.16 32.72 11.22 ;
			RECT 32 2.16 32.72 2.8 ;

		END 

		ANTENNADIFFAREA 3.828 LAYER MTL1  ;
	END Q
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 33.12 13.68 ;
			RECT 30.24 8.58 30.88 13.68 ;
			RECT 28.36 10.7 29 13.68 ;
			RECT 21.44 8.58 22.08 13.68 ;
			RECT 18.48 9.92 19.12 13.68 ;
			RECT 12.4 10.7 13.04 13.68 ;
			RECT 7.12 10.7 7.76 13.68 ;
			RECT 2.32 10.58 2.96 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 33.12 1.46 ;
			RECT 30.6 -0.48 31.24 2.76 ;
			RECT 26.28 -0.48 26.92 3.7 ;
			RECT 21.48 -0.48 22.12 3.44 ;
			RECT 17.96 -0.48 18.6 2.06 ;
			RECT 12.8 -0.48 13.44 2.78 ;
			RECT 7.74 -0.48 8.4 2.26 ;
			RECT 1.86 -0.48 2.5 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1.86 3.14 5.38 3.62 ;
			RECT 1.86 3.14 2.5 3.9 ;
			RECT 4.74 3.14 5.38 4.78 ;
			RECT 4.9 7.54 5.88 9.18 ;
			RECT 4.9 3.14 5.38 10.06 ;
			RECT 0.88 9.58 5.38 10.06 ;
			RECT 0.88 9.58 1.52 11.22 ;
			RECT 5.1 1.98 7.12 2.62 ;
			RECT 6.6 1.98 7.12 3.26 ;
			RECT 6.6 2.78 9.16 3.26 ;
			RECT 8.52 2.78 9.16 3.7 ;
			RECT 6.12 9.7 9.2 10.18 ;
			RECT 8.56 9.7 9.2 10.86 ;
			RECT 6.12 9.7 6.6 11.06 ;
			RECT 4.72 10.58 6.6 11.06 ;
			RECT 4.72 10.58 5.36 11.22 ;
			RECT 10.8 4.58 11.44 9.18 ;
			RECT 8.52 8.54 11.44 9.18 ;
			RECT 10.16 2.26 10.8 2.9 ;
			RECT 10.28 2.26 10.8 3.78 ;
			RECT 10.28 3.3 13.92 3.78 ;
			RECT 13.12 3.3 13.92 4.02 ;
			RECT 12.48 9.22 13.6 9.86 ;
			RECT 13.12 3.3 13.6 9.86 ;
			RECT 10.12 9.7 12.96 10.18 ;
			RECT 10.12 9.7 10.6 11.22 ;
			RECT 9.96 10.58 10.6 11.22 ;
			RECT 14.44 2.38 15.08 5.22 ;
			RECT 14.44 3.58 15.44 5.22 ;
			RECT 14.44 8.22 15.12 9.86 ;
			RECT 14.44 2.38 14.92 11.22 ;
			RECT 13.84 10.58 14.92 11.22 ;
			RECT 16.44 1.98 17.08 3.06 ;
			RECT 15.96 2.58 18.64 3.06 ;
			RECT 18.16 2.58 18.64 3.78 ;
			RECT 18.16 3.14 19.96 3.78 ;
			RECT 15.96 2.58 16.44 10.56 ;
			RECT 15.96 6.98 16.6 10.56 ;
			RECT 15.96 9.92 17.72 10.56 ;
			RECT 19.72 1.98 20.96 2.62 ;
			RECT 20.48 1.98 20.96 6.22 ;
			RECT 19.92 5.58 21.58 6.22 ;
			RECT 19.92 5.58 20.56 10.12 ;
			RECT 22.88 2.8 23.52 11.22 ;
			RECT 27.72 8.54 29.36 9.18 ;
			RECT 27.72 8.54 28.36 10.18 ;
			RECT 27.72 1.98 29.56 2.62 ;
			RECT 27.72 1.98 28.36 6.58 ;
			RECT 28.92 3.44 31.56 4.08 ;
			RECT 28.92 3.44 29.4 8.02 ;
			RECT 24.28 7.38 31.4 8.02 ;
			RECT 24.28 2.8 24.92 11.22 ;
			RECT 24.28 10.58 26.36 11.22 ;

	END

END DFMH

MACRO DFCSLQ
	CLASS CORE ;
	FOREIGN DFCSLQ 0 0  ;
	ORIGIN 0 0 ;
	SIZE 43.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN C
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER MTL1 ;
			RECT 32.6 6.28 33.24 9.04 ;
			RECT 30.64 6.28 33.24 6.92 ;
			RECT 30.64 4.96 32.04 6.92 ;
			RECT 31.4 3.54 32.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.821 LAYER MTL1  ;
	END C
	PIN D0
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 2.16 3.78 3.8 4.42 ;
			RECT 1.84 7.6 3.48 8.24 ;
			RECT 3 3.78 3.48 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.749 LAYER MTL1  ;
	END D0
	PIN D1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 5.28 8.24 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.749 LAYER MTL1  ;
	END D1
	PIN S1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.397 LAYER MTL1  ;
	END S1
	PIN SCIN
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 13.2 6.74 14 8.42 ;
			RECT 13.36 3.14 14 8.42 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.691 LAYER MTL1  ;
	END SCIN
	PIN SCEN
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 9.04 7.6 10.68 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.656 LAYER MTL1  ;
	END SCEN
	PIN SB
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 23.16 9.22 24.8 9.86 ;
			RECT 23.44 3.14 24.16 4.78 ;
			RECT 23.44 3.14 24.08 9.86 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.57 LAYER MTL1  ;
	END SB
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 42.16 1.98 42.8 11.22 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END Q
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 43.2 13.68 ;
			RECT 40.76 9.26 41.4 13.68 ;
			RECT 39.32 10.58 39.96 13.68 ;
			RECT 33.52 10.68 34.16 13.68 ;
			RECT 28.24 10.32 28.88 13.68 ;
			RECT 25.16 10.58 25.8 13.68 ;
			RECT 22.56 10.58 23.2 13.68 ;
			RECT 19.76 10.7 20.4 13.68 ;
			RECT 13.24 10.94 13.88 13.68 ;
			RECT 9.44 11.66 10.08 13.68 ;
			RECT 1 10.9 1.64 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 43.2 1.46 ;
			RECT 40.76 -0.48 41.4 2.66 ;
			RECT 35.22 -0.48 35.86 1.8 ;
			RECT 30.4 -0.48 31.04 2.54 ;
			RECT 24.16 -0.48 24.8 2.62 ;
			RECT 20.08 -0.48 20.72 2.62 ;
			RECT 13.16 -0.48 13.8 1.62 ;
			RECT 9.56 -0.48 10.2 2.26 ;
			RECT 1 -0.48 1.64 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1 2.78 5.04 3.26 ;
			RECT 1 2.78 1.64 3.9 ;
			RECT 4.44 2.78 5.04 5.62 ;
			RECT 4.44 3.98 5.56 5.62 ;
			RECT 4.44 7.94 6.66 8.58 ;
			RECT 4.44 2.78 4.92 10.2 ;
			RECT 1 9.54 4.92 10.2 ;
			RECT 11.72 3.14 12.36 4.42 ;
			RECT 8.72 3.78 12.36 4.42 ;
			RECT 11.2 3.78 11.68 10.14 ;
			RECT 14.56 8.06 15.2 9.42 ;
			RECT 11.2 8.94 15.2 9.42 ;
			RECT 11.2 8.94 11.72 10.14 ;
			RECT 11.08 9.5 11.72 10.14 ;
			RECT 12.24 9.94 15.24 10.42 ;
			RECT 14.76 9.94 15.24 11.22 ;
			RECT 5.48 9.4 6.12 11.14 ;
			RECT 12.24 9.94 12.72 11.14 ;
			RECT 5.48 10.66 12.72 11.14 ;
			RECT 14.76 10.58 16.44 11.22 ;
			RECT 15.8 1.98 16.44 2.62 ;
			RECT 10.72 2.14 16.44 2.62 ;
			RECT 10.72 2.14 11.2 3.26 ;
			RECT 5.56 2.78 11.2 3.26 ;
			RECT 5.56 2.78 6.2 3.46 ;
			RECT 17.8 3.14 18.44 4.78 ;
			RECT 17.8 3.14 18.28 9.06 ;
			RECT 16.68 7.42 18.28 9.06 ;
			RECT 17.44 1.98 18.08 2.62 ;
			RECT 17.44 2.14 19.48 2.62 ;
			RECT 19 3.14 21.08 3.8 ;
			RECT 19 9.22 20.76 9.86 ;
			RECT 19 2.14 19.48 10.18 ;
			RECT 17.2 9.7 19.48 10.18 ;
			RECT 17.2 9.7 17.84 11.22 ;
			RECT 21.52 1.98 22.16 2.62 ;
			RECT 21.6 1.98 22.08 5 ;
			RECT 20 4.52 21.76 5.16 ;
			RECT 21.28 4.52 21.76 11.22 ;
			RECT 20.28 7.86 21.92 8.5 ;
			RECT 21.28 7.86 21.92 11.22 ;
			RECT 21.16 10.58 21.92 11.22 ;
			RECT 25.98 1.98 27.2 2.62 ;
			RECT 25.98 1.98 26.46 4.78 ;
			RECT 26.32 4.3 27.22 6.18 ;
			RECT 26.32 4.3 26.8 10.7 ;
			RECT 26.32 10.06 27.44 10.7 ;
			RECT 28.76 3.54 30.54 4.18 ;
			RECT 28.76 3.54 29.24 8.54 ;
			RECT 28.76 7.9 29.4 8.54 ;
			RECT 27.76 1.98 28.64 2.62 ;
			RECT 27 3.14 28.24 3.78 ;
			RECT 30.64 8.26 31.76 8.9 ;
			RECT 27.76 1.98 28.24 9.54 ;
			RECT 27.32 8.9 28.24 9.54 ;
			RECT 27.32 9.06 31.28 9.54 ;
			RECT 30.64 8.26 31.28 11.22 ;
			RECT 31.92 1.98 33.06 2.62 ;
			RECT 32.58 1.98 33.06 3.96 ;
			RECT 32.58 3.32 34.28 3.96 ;
			RECT 33.8 8.4 34.6 9.06 ;
			RECT 33.8 3.32 34.28 10.04 ;
			RECT 32.08 9.56 34.28 10.04 ;
			RECT 32.08 9.56 32.76 11.22 ;
			RECT 33.58 1.98 34.22 2.8 ;
			RECT 33.58 2.32 35.28 2.8 ;
			RECT 34.8 2.32 35.28 5.18 ;
			RECT 35.12 9.42 37.64 10.06 ;
			RECT 35.12 4.54 35.6 11.22 ;
			RECT 34.92 10.58 35.6 11.22 ;
			RECT 37.88 1.98 38.52 2.8 ;
			RECT 36.12 2.32 38.52 2.8 ;
			RECT 36.12 2.32 36.76 8.9 ;
			RECT 36.12 8.42 38.76 8.9 ;
			RECT 38.28 8.42 38.76 11.22 ;
			RECT 36.36 10.58 38.76 11.22 ;
			RECT 37.28 3.32 40.56 3.8 ;
			RECT 39.92 3.32 40.56 4.3 ;
			RECT 37.28 3.32 37.76 7.5 ;
			RECT 37.28 7.02 40 7.5 ;
			RECT 39.28 7.02 40 9.74 ;

	END

END DFCSLQ

MACRO DFCRLSLQ
	CLASS CORE ;
	FOREIGN DFCRLSLQ 0 0  ;
	ORIGIN 0 0 ;
	SIZE 48.96 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN C
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER MTL1 ;
			RECT 38.36 6.28 39 9.04 ;
			RECT 36.4 7.6 39 8.24 ;
			RECT 36.82 6.28 39 8.24 ;
			RECT 36.82 3.76 37.46 8.24 ;
			RECT 36.4 6.28 39 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.821 LAYER MTL1  ;
	END C
	PIN D0
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 2.24 3.78 3.88 4.42 ;
			RECT 1.84 7.6 3.48 8.24 ;
			RECT 3 3.78 3.48 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.749 LAYER MTL1  ;
	END D0
	PIN D1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 5.26 8.24 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.749 LAYER MTL1  ;
	END D1
	PIN S1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.397 LAYER MTL1  ;
	END S1
	PIN SCIN
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 13.2 6.78 14 8.42 ;
			RECT 13.36 3.14 14 8.42 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.706 LAYER MTL1  ;
	END SCIN
	PIN SCEN
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 9 7.6 10.68 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.728 LAYER MTL1  ;
	END SCEN
	PIN RB
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 26.48 4.54 27.16 5.18 ;
			RECT 25.54 6.28 26.96 8.24 ;
			RECT 26.48 4.54 26.96 8.24 ;
			RECT 25.54 6.28 26.36 9.56 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.562 LAYER MTL1  ;
	END RB
	PIN SB
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 28.72 8.9 30.4 9.54 ;
			RECT 29.92 5.54 30.4 9.54 ;
			RECT 28.68 5.54 30.4 6.18 ;
			RECT 19 3.14 21.08 3.8 ;
			RECT 19 9.46 20.76 10.14 ;
			RECT 19 7.6 19.76 10.14 ;
			RECT 19 6.28 19.76 6.92 ;
			RECT 19 3.14 19.48 10.14 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.872 LAYER MTL1  ;
	END SB
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 47.92 1.98 48.56 11.22 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END Q
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 48.96 13.68 ;
			RECT 46.52 9.12 47.16 13.68 ;
			RECT 45.08 10.58 45.72 13.68 ;
			RECT 39.28 10.68 39.92 13.68 ;
			RECT 34 10.32 34.64 13.68 ;
			RECT 29.64 11.06 30.28 13.68 ;
			RECT 24.72 10.58 25.36 13.68 ;
			RECT 19.76 11.66 20.4 13.68 ;
			RECT 13.24 10.94 13.88 13.68 ;
			RECT 9.44 11.66 10.08 13.68 ;
			RECT 1 10.9 1.64 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 48.96 1.46 ;
			RECT 46.52 -0.48 47.16 2.66 ;
			RECT 40.98 -0.48 41.62 1.8 ;
			RECT 35.96 -0.48 36.6 2.54 ;
			RECT 27.8 -0.48 28.44 2.5 ;
			RECT 20.08 -0.48 20.72 2.58 ;
			RECT 13.16 -0.48 13.8 1.62 ;
			RECT 9.56 -0.48 10.2 2.26 ;
			RECT 1 -0.48 1.64 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1 2.78 5.04 3.26 ;
			RECT 1 2.78 1.64 3.9 ;
			RECT 4.44 2.78 5.04 5.62 ;
			RECT 4.44 3.98 5.56 5.62 ;
			RECT 4.44 7.94 6.66 8.58 ;
			RECT 4.44 2.78 4.92 10.2 ;
			RECT 1 9.54 4.92 10.2 ;
			RECT 11.72 3.14 12.36 4.42 ;
			RECT 8.72 3.78 12.36 4.42 ;
			RECT 11.2 3.78 11.68 10.14 ;
			RECT 14.56 8.06 15.2 9.42 ;
			RECT 11.2 8.94 15.2 9.42 ;
			RECT 11.2 8.94 11.72 10.14 ;
			RECT 11.08 9.5 11.72 10.14 ;
			RECT 12.24 9.94 15.24 10.42 ;
			RECT 14.76 9.94 15.24 11.22 ;
			RECT 5.48 9.4 6.12 11.14 ;
			RECT 12.24 9.94 12.72 11.14 ;
			RECT 5.48 10.66 12.72 11.14 ;
			RECT 14.76 10.58 16.44 11.22 ;
			RECT 15.8 1.98 16.44 2.62 ;
			RECT 10.72 2.14 16.44 2.62 ;
			RECT 10.72 2.14 11.2 3.26 ;
			RECT 5.56 2.78 11.2 3.26 ;
			RECT 5.56 2.78 6.2 3.46 ;
			RECT 16.96 4.8 18.44 5.44 ;
			RECT 16.96 4.8 17.44 9.06 ;
			RECT 16.76 7.42 17.44 9.06 ;
			RECT 23 2.98 23.64 5 ;
			RECT 20 4.52 23.64 5 ;
			RECT 20 4.52 21.96 5.16 ;
			RECT 21.48 4.52 21.96 8.54 ;
			RECT 21.68 7.9 22.32 10.14 ;
			RECT 17.44 1.98 18.08 3.62 ;
			RECT 15.76 3.14 18.08 3.62 ;
			RECT 24.16 3.14 24.8 3.78 ;
			RECT 15.76 3.14 16.24 10.06 ;
			RECT 24.16 3.14 24.64 9.7 ;
			RECT 22.84 9.06 24.64 9.7 ;
			RECT 15.76 9.58 17.84 10.06 ;
			RECT 22.84 9.06 23.32 11.14 ;
			RECT 17.2 10.66 23.32 11.14 ;
			RECT 17.2 9.58 17.84 11.22 ;
			RECT 21.48 1.98 25.16 2.46 ;
			RECT 21.48 1.98 22.12 2.62 ;
			RECT 24.52 1.98 25.16 2.62 ;
			RECT 26.16 1.98 26.8 4.02 ;
			RECT 25.32 3.54 30.2 4.02 ;
			RECT 29.72 3.54 30.2 4.78 ;
			RECT 29.72 4.14 30.36 4.78 ;
			RECT 25.32 3.54 25.8 5.18 ;
			RECT 25.16 4.54 25.8 5.18 ;
			RECT 27.68 3.54 28.16 9.54 ;
			RECT 26.88 8.9 28.16 9.54 ;
			RECT 26.88 8.9 27.4 11.22 ;
			RECT 26.28 10.58 27.4 11.22 ;
			RECT 30.72 2.98 31.4 3.62 ;
			RECT 30.92 5.54 32.68 6.18 ;
			RECT 30.92 2.98 31.4 10.54 ;
			RECT 28.12 10.06 32.68 10.54 ;
			RECT 28.12 10.06 28.76 11.22 ;
			RECT 32.04 10.06 32.68 11.22 ;
			RECT 29.2 1.98 32.76 2.46 ;
			RECT 29.2 1.98 29.84 2.62 ;
			RECT 32.12 1.98 32.76 3.34 ;
			RECT 34.4 3.76 36.1 4.4 ;
			RECT 34.4 3.76 34.88 8.54 ;
			RECT 34.4 7.9 35.04 8.54 ;
			RECT 33.4 1.98 34.2 2.62 ;
			RECT 31.92 4.18 33.88 4.82 ;
			RECT 33.4 1.98 33.88 9.54 ;
			RECT 33.04 8.9 33.88 9.54 ;
			RECT 36.44 8.9 37.56 9.54 ;
			RECT 33.04 9.06 37.56 9.54 ;
			RECT 36.4 9.06 37.04 11.22 ;
			RECT 37.6 1.98 38.46 2.62 ;
			RECT 37.98 1.98 38.46 4.62 ;
			RECT 37.98 4.14 40.98 4.62 ;
			RECT 40.34 3.36 40.98 5 ;
			RECT 40 8.4 40.8 9.06 ;
			RECT 40 4.14 40.48 10.04 ;
			RECT 38.08 9.56 40.48 10.04 ;
			RECT 38.08 9.56 38.56 11.22 ;
			RECT 37.84 10.5 38.56 11.22 ;
			RECT 38.98 1.98 39.98 2.8 ;
			RECT 38.98 2.32 41.98 2.8 ;
			RECT 38.98 1.98 39.62 3.62 ;
			RECT 41.5 2.32 41.98 10.06 ;
			RECT 41.5 9.42 43.4 10.06 ;
			RECT 41.12 9.58 41.6 11.22 ;
			RECT 40.68 10.58 41.6 11.22 ;
			RECT 42.5 1.98 44.28 2.62 ;
			RECT 42.5 1.98 43.14 8.9 ;
			RECT 42.5 8.42 44.52 8.9 ;
			RECT 44.04 8.42 44.52 11.22 ;
			RECT 42.12 10.58 44.52 11.22 ;
			RECT 43.66 3.66 46.32 4.3 ;
			RECT 43.66 3.66 44.14 7.5 ;
			RECT 43.66 7.02 45.76 7.5 ;
			RECT 45.04 7.02 45.76 9.74 ;

	END

END DFCRLSLQ

MACRO DFCRLQ
	CLASS CORE ;
	FOREIGN DFCRLQ 0 0  ;
	ORIGIN 0 0 ;
	SIZE 47.52 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN C
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER MTL1 ;
			RECT 36.92 6.28 37.6 9.04 ;
			RECT 34.96 7.6 37.6 8.24 ;
			RECT 35.38 6.28 37.6 8.24 ;
			RECT 35.38 3.76 36.02 8.24 ;
			RECT 34.96 6.28 37.6 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.821 LAYER MTL1  ;
	END C
	PIN D0
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 2.16 3.78 3.8 4.42 ;
			RECT 1.84 7.6 3.48 8.24 ;
			RECT 3 3.78 3.48 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.792 LAYER MTL1  ;
	END D0
	PIN D1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 5.28 8.24 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.792 LAYER MTL1  ;
	END D1
	PIN S1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.44 LAYER MTL1  ;
	END S1
	PIN SCIN
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 13.2 6.78 14 8.42 ;
			RECT 13.36 3.14 14 8.42 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.706 LAYER MTL1  ;
	END SCIN
	PIN SCEN
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 9.04 7.6 10.68 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.728 LAYER MTL1  ;
	END SCEN
	PIN RB
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 26.76 8.9 28.4 9.56 ;
			RECT 27.76 3.14 28.4 9.56 ;
			RECT 27.24 3.14 28.4 4.78 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.562 LAYER MTL1  ;
	END RB
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 46.48 1.98 47.12 11.22 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END Q
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 47.52 13.68 ;
			RECT 45.08 9.1 45.72 13.68 ;
			RECT 43.64 10.58 44.28 13.68 ;
			RECT 37.84 10.68 38.48 13.68 ;
			RECT 32.56 10.74 33.2 13.68 ;
			RECT 27.96 10.38 28.6 13.68 ;
			RECT 24.04 11.22 24.68 13.68 ;
			RECT 20.2 10.7 20.84 13.68 ;
			RECT 13.24 10.94 13.88 13.68 ;
			RECT 9.44 11.66 10.08 13.68 ;
			RECT 1 10.9 1.64 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 47.52 1.46 ;
			RECT 45.08 -0.48 45.72 2.66 ;
			RECT 39.54 -0.48 40.18 1.8 ;
			RECT 34.52 -0.48 35.16 2.82 ;
			RECT 30.66 -0.48 31.32 2.62 ;
			RECT 27.88 -0.48 28.52 2.62 ;
			RECT 24.8 -0.48 25.44 2.14 ;
			RECT 21.52 -0.48 22.16 1.78 ;
			RECT 14.58 -0.48 15.22 1.62 ;
			RECT 9.56 -0.48 10.2 2.26 ;
			RECT 1 -0.48 1.64 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1 2.78 5.04 3.26 ;
			RECT 1 2.78 1.64 3.9 ;
			RECT 4.44 2.78 5.04 5.62 ;
			RECT 4.44 3.98 5.56 5.62 ;
			RECT 4.44 7.82 6.66 8.46 ;
			RECT 4.44 2.78 4.92 10.2 ;
			RECT 1 9.54 4.92 10.2 ;
			RECT 11.72 3.14 12.36 4.42 ;
			RECT 8.72 3.78 12.36 4.42 ;
			RECT 11.2 3.78 11.68 10.14 ;
			RECT 14.56 8.06 15.2 9.42 ;
			RECT 11.2 8.94 15.2 9.42 ;
			RECT 11.2 8.94 11.72 10.14 ;
			RECT 11.08 9.5 11.72 10.14 ;
			RECT 12.24 9.94 15.24 10.42 ;
			RECT 14.76 9.94 15.24 11.22 ;
			RECT 5.48 9.4 6.12 11.14 ;
			RECT 12.24 9.94 12.72 11.14 ;
			RECT 5.48 10.66 12.72 11.14 ;
			RECT 14.76 10.58 16.44 11.22 ;
			RECT 17.22 1.98 17.86 2.62 ;
			RECT 10.72 2.14 17.86 2.62 ;
			RECT 10.72 2.14 11.2 3.26 ;
			RECT 5.56 2.78 11.2 3.26 ;
			RECT 5.56 2.78 6.2 3.46 ;
			RECT 19.48 3.3 20.12 9.06 ;
			RECT 16.32 8.42 20.12 9.06 ;
			RECT 23.16 1.98 23.8 2.78 ;
			RECT 21.8 2.3 23.8 2.78 ;
			RECT 21.8 2.3 22.44 8.34 ;
			RECT 23.96 7.7 24.6 10.7 ;
			RECT 21.64 10.22 24.6 10.7 ;
			RECT 21.64 10.22 22.34 10.86 ;
			RECT 18.86 1.98 19.54 2.78 ;
			RECT 18.86 2.3 21.12 2.78 ;
			RECT 24.32 2.66 24.96 3.78 ;
			RECT 22.96 3.3 24.96 3.78 ;
			RECT 20.64 9.06 23.44 9.7 ;
			RECT 22.96 3.3 23.44 9.7 ;
			RECT 20.64 2.3 21.12 10.18 ;
			RECT 17.76 9.7 21.12 10.18 ;
			RECT 17.76 9.7 18.4 11.22 ;
			RECT 25.96 1.98 26.88 2.62 ;
			RECT 25.96 1.98 26.44 4.94 ;
			RECT 24.12 4.3 26.44 4.94 ;
			RECT 25.12 4.3 25.6 10.7 ;
			RECT 25.56 10.22 27.2 11.22 ;
			RECT 29.28 1.98 30.14 2.62 ;
			RECT 29.66 1.98 30.14 3.62 ;
			RECT 29.66 3.14 30.92 3.62 ;
			RECT 30.28 3.14 30.92 5.4 ;
			RECT 30.36 3.14 30.92 11.22 ;
			RECT 30.36 9.44 31 11.22 ;
			RECT 32.84 3.76 34.66 4.4 ;
			RECT 32.84 3.76 33.32 8.38 ;
			RECT 32.6 7.7 33.32 8.38 ;
			RECT 31.84 1.98 32.76 2.62 ;
			RECT 31.84 1.98 32.32 4.38 ;
			RECT 34.96 8.9 36.12 9.54 ;
			RECT 31.56 3.74 32.04 10.22 ;
			RECT 31.56 9.56 35.6 10.22 ;
			RECT 34.96 8.9 35.6 11.22 ;
			RECT 36.16 1.98 37.02 2.62 ;
			RECT 36.54 1.98 37.02 4.62 ;
			RECT 38.9 3.36 39.54 4.62 ;
			RECT 36.54 4.14 39.54 4.62 ;
			RECT 38.56 7.42 39.36 9.06 ;
			RECT 38.56 4.14 39.04 10.04 ;
			RECT 36.64 9.56 39.04 10.04 ;
			RECT 36.64 9.56 37.12 11.22 ;
			RECT 36.4 10.5 37.12 11.22 ;
			RECT 37.54 1.98 38.54 2.8 ;
			RECT 37.54 2.32 40.54 2.8 ;
			RECT 37.54 1.98 38.18 3.62 ;
			RECT 40.06 2.32 40.54 10.06 ;
			RECT 40.06 8.9 40.76 10.06 ;
			RECT 39.56 9.58 40.76 10.06 ;
			RECT 39.56 9.58 40.04 11.22 ;
			RECT 39.24 10.58 40.04 11.22 ;
			RECT 41.28 1.98 42.84 2.62 ;
			RECT 41.06 6.5 41.76 8.18 ;
			RECT 41.28 1.98 41.76 11.22 ;
			RECT 40.68 10.58 41.76 11.22 ;
			RECT 42.32 3.66 44.88 4.3 ;
			RECT 42.32 3.66 42.8 7.6 ;
			RECT 42.32 7.02 44.32 7.6 ;
			RECT 43.54 7.02 44.32 9.74 ;

	END

END DFCRLQ

MACRO DFCQ
	CLASS CORE ;
	FOREIGN DFCQ 0 0  ;
	ORIGIN 0 0 ;
	SIZE 40.32 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN C
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER MTL1 ;
			RECT 29.2 7.6 31.28 8.24 ;
			RECT 29.62 6.28 31.28 8.24 ;
			RECT 30.44 6.28 31.08 9.04 ;
			RECT 29.62 3.76 30.26 8.24 ;
			RECT 29.2 6.28 31.28 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.821 LAYER MTL1  ;
	END C
	PIN D0
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 2.16 3.78 3.84 4.42 ;
			RECT 1.84 7.6 3.48 8.24 ;
			RECT 3 3.78 3.48 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.706 LAYER MTL1  ;
	END D0
	PIN D1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 5.28 8.24 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.706 LAYER MTL1  ;
	END D1
	PIN S1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.354 LAYER MTL1  ;
	END S1
	PIN SCIN
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 13.2 6.78 14 8.42 ;
			RECT 13.36 3.14 14 8.42 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.648 LAYER MTL1  ;
	END SCIN
	PIN SCEN
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 9.02 7.6 10.66 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.656 LAYER MTL1  ;
	END SCEN
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 39.28 1.98 39.92 11.22 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END Q
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 40.32 13.68 ;
			RECT 36.48 10.58 38.52 13.68 ;
			RECT 37.88 9.1 38.52 13.68 ;
			RECT 31 10.68 31.64 13.68 ;
			RECT 25.72 10.14 26.36 13.68 ;
			RECT 22.68 10.38 23.32 13.68 ;
			RECT 19.64 10.7 20.28 13.68 ;
			RECT 13.24 10.94 13.88 13.68 ;
			RECT 9.44 11.66 10.08 13.68 ;
			RECT 1 10.9 1.64 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 40.32 1.46 ;
			RECT 37.88 -0.48 38.52 2.26 ;
			RECT 33.78 -0.48 34.42 1.8 ;
			RECT 28.76 -0.48 29.4 2.82 ;
			RECT 23.26 -0.48 23.9 2.14 ;
			RECT 20.18 -0.48 20.82 1.78 ;
			RECT 13.16 -0.48 13.8 1.62 ;
			RECT 9.56 -0.48 10.2 2.26 ;
			RECT 1 -0.48 1.64 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1 2.78 5.04 3.26 ;
			RECT 1 2.78 1.64 3.9 ;
			RECT 4.44 2.78 5.04 5.62 ;
			RECT 4.44 3.98 5.56 5.62 ;
			RECT 4.44 8.06 6.66 8.7 ;
			RECT 4.44 2.78 4.92 10.2 ;
			RECT 1 9.54 4.92 10.2 ;
			RECT 11.72 3.14 12.36 4.42 ;
			RECT 8.72 3.78 12.36 4.42 ;
			RECT 11.2 3.78 11.68 10.14 ;
			RECT 14.56 8.06 15.2 9.42 ;
			RECT 11.2 8.94 15.2 9.42 ;
			RECT 11.2 8.94 11.72 10.14 ;
			RECT 11.08 9.5 11.72 10.14 ;
			RECT 12.24 9.94 15.24 10.42 ;
			RECT 14.76 9.94 15.24 11.22 ;
			RECT 5.48 9.4 6.12 11.14 ;
			RECT 12.24 9.94 12.72 11.14 ;
			RECT 5.48 10.66 12.72 11.14 ;
			RECT 14.76 10.58 16.44 11.22 ;
			RECT 15.8 1.98 16.44 2.62 ;
			RECT 10.72 2.14 16.44 2.62 ;
			RECT 10.72 2.14 11.2 3.26 ;
			RECT 5.56 2.78 11.2 3.26 ;
			RECT 5.56 2.78 6.2 3.46 ;
			RECT 17.88 3.3 18.52 7.9 ;
			RECT 16.68 7.42 18.52 7.9 ;
			RECT 16.68 7.42 17.32 9.06 ;
			RECT 17.52 1.98 18.2 2.78 ;
			RECT 17.52 2.3 19.62 2.78 ;
			RECT 19.14 4.04 20.18 5.68 ;
			RECT 19.14 2.3 19.62 10.18 ;
			RECT 17.2 9.7 19.62 10.18 ;
			RECT 17.2 9.7 17.84 11.22 ;
			RECT 21.62 1.98 22.26 3.32 ;
			RECT 20.14 2.68 22.26 3.32 ;
			RECT 20.7 2.68 21.34 9.62 ;
			RECT 20.8 2.68 21.34 11.22 ;
			RECT 20.8 10.56 21.92 11.22 ;
			RECT 22.16 4.04 22.84 9.7 ;
			RECT 24.9 1.98 25.56 3.24 ;
			RECT 24.08 2.76 25.56 3.24 ;
			RECT 24.08 2.76 24.72 11.22 ;
			RECT 27.08 3.76 28.9 4.4 ;
			RECT 27.08 3.76 27.56 8.26 ;
			RECT 26.24 7.62 27.56 8.26 ;
			RECT 26.08 1.98 27 2.62 ;
			RECT 26.08 1.98 26.56 4.4 ;
			RECT 25.24 3.76 26.56 4.4 ;
			RECT 25.24 3.76 25.72 9.62 ;
			RECT 25.24 8.98 29.24 9.62 ;
			RECT 28.12 8.98 28.76 11.22 ;
			RECT 30.4 1.98 31.26 2.62 ;
			RECT 30.78 1.98 31.26 4.62 ;
			RECT 33.14 3.36 33.78 4.62 ;
			RECT 30.78 4.14 33.78 4.62 ;
			RECT 31.84 7.42 32.52 9.06 ;
			RECT 31.84 4.14 32.32 10.04 ;
			RECT 30 9.56 32.32 10.04 ;
			RECT 30 9.56 30.48 11.22 ;
			RECT 29.56 10.5 30.48 11.22 ;
			RECT 31.78 1.98 32.78 2.8 ;
			RECT 31.78 2.32 34.78 2.8 ;
			RECT 31.78 1.98 32.42 3.62 ;
			RECT 34.3 2.32 34.78 5.62 ;
			RECT 33.28 5.14 34.78 5.62 ;
			RECT 33.28 5.14 33.76 10.06 ;
			RECT 33.28 9.42 34.96 10.06 ;
			RECT 32.84 9.58 33.32 11.22 ;
			RECT 32.4 10.56 33.32 11.22 ;
			RECT 35.48 1.98 37.08 2.62 ;
			RECT 35.48 1.98 36 6.82 ;
			RECT 35.48 5.18 37.28 6.82 ;
			RECT 34.28 7.06 35.96 8.7 ;
			RECT 35.48 1.98 35.96 11.22 ;
			RECT 33.84 10.58 35.96 11.22 ;

	END

END DFCQ

MACRO DFCHSL
	CLASS CORE ;
	FOREIGN DFCHSL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 43.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN C
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER MTL1 ;
			RECT 29.08 3.14 29.84 8.72 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.821 LAYER MTL1  ;
	END C
	PIN D0
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 2.16 3.78 3.8 4.42 ;
			RECT 1.84 7.6 3.48 8.24 ;
			RECT 3 3.78 3.48 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.763 LAYER MTL1  ;
	END D0
	PIN D1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 5.28 8.24 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.763 LAYER MTL1  ;
	END D1
	PIN S1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.411 LAYER MTL1  ;
	END S1
	PIN SCIN
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 13.2 6.74 14 8.42 ;
			RECT 13.36 3.14 14 8.42 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.734 LAYER MTL1  ;
	END SCIN
	PIN SCEN
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 9.04 7.6 10.68 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.915 LAYER MTL1  ;
	END SCEN
	PIN SB
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 23.44 3.74 24.16 4.38 ;
			RECT 22.28 8.78 24.08 9.42 ;
			RECT 23.44 3.64 24.08 9.42 ;
			RECT 22.28 8.78 22.92 9.86 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.779 LAYER MTL1  ;
	END SB
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 40.24 7.6 42.8 8.26 ;
			RECT 42.16 2.2 42.8 8.26 ;
			RECT 40.24 7.6 40.88 11.04 ;

		END 

		ANTENNADIFFAREA 4.598 LAYER MTL1  ;
	END Q
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 43.2 13.68 ;
			RECT 41.64 8.88 42.28 13.68 ;
			RECT 38.84 8.24 39.48 13.68 ;
			RECT 35.56 10.7 36.2 13.68 ;
			RECT 29.96 10.24 30.6 13.68 ;
			RECT 22.66 10.58 23.3 13.68 ;
			RECT 19.76 10.7 20.4 13.68 ;
			RECT 13.24 10.94 13.88 13.68 ;
			RECT 9.44 11.66 10.08 13.68 ;
			RECT 1 10.9 1.64 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 43.2 1.46 ;
			RECT 39.76 -0.48 40.4 2.84 ;
			RECT 34.48 -0.48 35.12 2.78 ;
			RECT 28.6 -0.48 29.24 2.5 ;
			RECT 24.16 -0.48 24.8 2.62 ;
			RECT 20.08 -0.48 20.72 2.62 ;
			RECT 13.16 -0.48 13.8 1.62 ;
			RECT 9.56 -0.48 10.2 2.26 ;
			RECT 1 -0.48 1.64 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1 2.78 5.04 3.26 ;
			RECT 1 2.78 1.64 3.9 ;
			RECT 4.44 2.78 5.04 5.62 ;
			RECT 4.44 3.98 5.56 5.62 ;
			RECT 4.44 7.86 6.66 8.5 ;
			RECT 4.44 2.78 4.92 10.2 ;
			RECT 1 9.54 4.92 10.2 ;
			RECT 11.72 3.14 12.36 4.42 ;
			RECT 8.72 3.78 12.36 4.42 ;
			RECT 11.2 3.78 11.68 10.14 ;
			RECT 14.56 6.9 15.2 9.42 ;
			RECT 11.2 8.94 15.2 9.42 ;
			RECT 11.2 8.94 11.72 10.14 ;
			RECT 11.08 9.5 11.72 10.14 ;
			RECT 12.24 9.94 15.24 10.42 ;
			RECT 14.76 9.94 15.24 11.22 ;
			RECT 5.48 9.4 6.12 11.14 ;
			RECT 12.24 9.94 12.72 11.14 ;
			RECT 5.48 10.66 12.72 11.14 ;
			RECT 14.76 10.58 16.44 11.22 ;
			RECT 15.8 1.98 16.44 2.62 ;
			RECT 10.72 2.14 16.44 2.62 ;
			RECT 10.72 2.14 11.2 3.26 ;
			RECT 5.56 2.78 11.2 3.26 ;
			RECT 5.56 2.78 6.2 3.46 ;
			RECT 17.8 3.14 18.44 4.78 ;
			RECT 17.8 3.14 18.28 9.18 ;
			RECT 16.68 7.54 18.28 9.18 ;
			RECT 17.44 1.98 18.08 2.62 ;
			RECT 17.44 2.14 19.48 2.62 ;
			RECT 19 3.14 21.08 3.8 ;
			RECT 19 9.22 20.76 9.86 ;
			RECT 19 2.14 19.48 10.18 ;
			RECT 17.2 9.7 19.48 10.18 ;
			RECT 17.2 9.7 17.84 11.22 ;
			RECT 21.52 1.98 22.16 2.62 ;
			RECT 21.6 1.98 22.08 5.22 ;
			RECT 20.12 4.74 21.76 5.38 ;
			RECT 20.12 7.78 21.76 8.42 ;
			RECT 21.28 4.74 21.76 11.22 ;
			RECT 21.16 10.58 21.8 11.22 ;
			RECT 25.56 1.98 26.2 8.06 ;
			RECT 24.6 7.44 26.2 8.06 ;
			RECT 24.6 7.44 25.24 11.22 ;
			RECT 26.96 1.98 27.6 9.22 ;
			RECT 26 8.58 27.6 9.22 ;
			RECT 26 8.58 26.64 11.22 ;
			RECT 30 1.98 31.12 2.62 ;
			RECT 30.4 1.98 31.12 8.46 ;
			RECT 30.4 6.82 31.24 8.46 ;
			RECT 30.4 1.98 30.96 9.72 ;
			RECT 28.56 9.24 30.96 9.72 ;
			RECT 28.56 9.24 29.24 10.8 ;
			RECT 31.84 2.1 33.48 2.76 ;
			RECT 31.84 2.1 33.2 3.76 ;
			RECT 32.56 2.1 33.2 10.06 ;
			RECT 31.48 9.42 33.2 10.06 ;
			RECT 37.12 1.98 37.76 2.78 ;
			RECT 35.78 2.28 37.76 2.78 ;
			RECT 35.78 2.28 36.26 4.9 ;
			RECT 35.12 4.26 36.26 4.9 ;
			RECT 35.48 6.94 36.12 8.58 ;
			RECT 35.48 7.94 37.84 8.58 ;
			RECT 37.2 7.94 37.84 11.14 ;
			RECT 37.12 3.46 38.4 4.1 ;
			RECT 37.76 3.46 38.4 6.34 ;
			RECT 33.76 5.7 41.52 6.34 ;
			RECT 40.88 4.84 41.52 6.5 ;
			RECT 33.76 5.7 34.56 7.5 ;
			RECT 33.76 5.7 34.24 11.22 ;
			RECT 32.92 10.58 34.24 11.22 ;

	END

END DFCHSL

MACRO DFCHRL
	CLASS CORE ;
	FOREIGN DFCHRL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 47.52 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN C
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER MTL1 ;
			RECT 29.04 4.46 30.68 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.821 LAYER MTL1  ;
	END C
	PIN D0
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 7.6 3.54 8.24 ;
			RECT 2.84 3.78 3.32 8.24 ;
			RECT 2.68 3.78 3.32 5.42 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.763 LAYER MTL1  ;
	END D0
	PIN D1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 6.28 7.52 6.92 ;
			RECT 6.88 5.28 7.52 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.763 LAYER MTL1  ;
	END D1
	PIN S1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.411 LAYER MTL1  ;
	END S1
	PIN SCIN
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 11.92 3.9 12.58 8.42 ;
			RECT 11.92 3.64 12.56 8.42 ;
			RECT 11.2 3.9 12.58 4.54 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.734 LAYER MTL1  ;
	END SCIN
	PIN SCEN
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 9.04 7.6 9.68 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.915 LAYER MTL1  ;
	END SCEN
	PIN RB
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 23.16 9.2 24.8 9.86 ;
			RECT 23.44 3.14 24.08 9.86 ;
			RECT 23 3.14 24.08 4.96 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.562 LAYER MTL1  ;
	END RB
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 46.44 2.1 47.14 11.14 ;
			RECT 43.78 3.82 47.14 4.46 ;

		END 

		ANTENNADIFFAREA 6.368 LAYER MTL1  ;
	END Q
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 47.52 13.68 ;
			RECT 42.3 8.4 42.94 13.68 ;
			RECT 39.84 10.9 40.48 13.68 ;
			RECT 32.72 10.42 33.36 13.68 ;
			RECT 29.12 9.56 29.76 13.68 ;
			RECT 22.12 11.42 22.76 13.68 ;
			RECT 17.08 11.32 17.72 13.68 ;
			RECT 9.16 10.94 10.96 13.68 ;
			RECT 1 10.9 1.64 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 47.52 1.46 ;
			RECT 44.04 -0.48 45.68 2.7 ;
			RECT 40.48 -0.48 41.18 1.6 ;
			RECT 37.8 -0.48 38.44 2.34 ;
			RECT 31.4 -0.48 32.04 2.94 ;
			RECT 27.68 -0.48 28.32 2.52 ;
			RECT 23.64 -0.48 24.28 2.62 ;
			RECT 20.56 -0.48 21.2 2.62 ;
			RECT 17.68 -0.48 18.32 2.62 ;
			RECT 9.32 -0.48 9.96 2.26 ;
			RECT 1 -0.48 1.64 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1 2.78 4.32 3.26 ;
			RECT 1 2.78 1.64 3.9 ;
			RECT 3.84 2.78 4.32 5.62 ;
			RECT 4.2 3.98 4.88 8.46 ;
			RECT 4.2 7.82 6.4 8.46 ;
			RECT 4.2 3.98 4.72 10.2 ;
			RECT 1 9.54 4.72 10.2 ;
			RECT 7.96 3.78 10.68 4.42 ;
			RECT 10.2 3.78 10.68 9.42 ;
			RECT 10.2 8.66 11.16 9.42 ;
			RECT 10.2 8.94 13.16 9.42 ;
			RECT 12.52 8.94 13.16 9.78 ;
			RECT 5.24 9.4 5.88 10.42 ;
			RECT 5.24 9.94 11.96 10.42 ;
			RECT 11.48 9.94 11.96 11.06 ;
			RECT 11.48 10.54 13.8 11.06 ;
			RECT 13.16 10.54 13.8 11.22 ;
			RECT 13.2 1.98 13.84 2.62 ;
			RECT 10.92 2.14 13.84 2.62 ;
			RECT 10.92 2.14 11.4 3.26 ;
			RECT 4.88 2.78 11.4 3.26 ;
			RECT 4.88 2.78 5.52 3.46 ;
			RECT 15.52 3.3 16.16 4.94 ;
			RECT 15.52 3.3 16 9.78 ;
			RECT 14.04 8.14 16 9.78 ;
			RECT 18.84 1.98 19.76 2.62 ;
			RECT 18.84 1.98 19.32 3.64 ;
			RECT 17.68 3.16 19.32 3.64 ;
			RECT 17.68 3.16 18.32 8.78 ;
			RECT 19.84 8.14 20.48 11.22 ;
			RECT 19.72 10.56 20.48 11.22 ;
			RECT 14.84 1.98 15.52 2.78 ;
			RECT 14.84 2.3 17.16 2.78 ;
			RECT 19.84 3.14 20.48 4.66 ;
			RECT 18.84 4.18 20.48 4.66 ;
			RECT 18.84 4.18 19.32 10.04 ;
			RECT 16.68 9.5 19.2 10.14 ;
			RECT 16.68 2.3 17.16 10.78 ;
			RECT 14.56 10.3 17.16 10.78 ;
			RECT 14.56 10.3 15.2 11.22 ;
			RECT 21.72 1.98 22.64 2.62 ;
			RECT 21.72 1.98 22.2 3.62 ;
			RECT 21 3.14 21.84 4.78 ;
			RECT 21 3.14 21.48 10.9 ;
			RECT 21 10.42 26.28 10.9 ;
			RECT 23.64 10.42 26.28 11.22 ;
			RECT 29.08 1.98 29.72 3.84 ;
			RECT 26.2 3.36 29.72 3.84 ;
			RECT 26.2 3.36 26.68 9.86 ;
			RECT 26.04 5.72 26.68 9.86 ;
			RECT 26.04 9.38 28.32 9.86 ;
			RECT 27.68 9.38 28.32 10.02 ;
			RECT 30.24 1.98 30.88 3.94 ;
			RECT 30.24 3.46 31.86 3.94 ;
			RECT 31.38 3.46 31.86 10.2 ;
			RECT 30.48 9.56 31.86 10.2 ;
			RECT 32.64 4.46 33.28 7.86 ;
			RECT 32.8 2.3 33.44 3.94 ;
			RECT 32.8 3.46 34.28 3.94 ;
			RECT 33.8 3.46 34.28 9.26 ;
			RECT 33.64 8.62 34.28 9.26 ;
			RECT 35.8 2.46 36.8 3.1 ;
			RECT 35.8 2.46 36.44 9.82 ;
			RECT 35.8 8.18 37.42 9.82 ;
			RECT 39.18 7.06 39.88 10.3 ;
			RECT 42.12 1.98 42.76 3.34 ;
			RECT 38.48 2.86 42.76 3.34 ;
			RECT 38.48 2.86 39.12 5.38 ;
			RECT 34.52 2.3 35.28 2.94 ;
			RECT 40.48 3.88 41.12 6.54 ;
			RECT 37.94 5.9 45.8 6.54 ;
			RECT 34.8 2.3 35.28 11.18 ;
			RECT 37.94 5.9 38.5 11.18 ;
			RECT 34.8 10.34 38.5 11.18 ;

	END

END DFCHRL

MACRO DFCH
	CLASS CORE ;
	FOREIGN DFCH 0 0  ;
	ORIGIN 0 0 ;
	SIZE 40.32 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN C
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER MTL1 ;
			RECT 24.88 8 26.54 8.64 ;
			RECT 24.88 4.96 25.52 8.64 ;
			RECT 24.16 4.96 25.52 5.6 ;
			RECT 24.16 3.58 24.8 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.821 LAYER MTL1  ;
	END C
	PIN D0
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 2.16 3.78 3.84 4.42 ;
			RECT 1.84 7.6 3.48 8.24 ;
			RECT 3 3.78 3.48 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.763 LAYER MTL1  ;
	END D0
	PIN D1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 5.28 8.24 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.763 LAYER MTL1  ;
	END D1
	PIN S1
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.411 LAYER MTL1  ;
	END S1
	PIN SCIN
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 13.36 6.78 14.52 8.42 ;
			RECT 13.36 3.14 14.44 4.82 ;
			RECT 13.36 3.14 14 8.42 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.691 LAYER MTL1  ;
	END SCIN
	PIN SCEN
		DIRECTION INPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 9.02 7.6 10.66 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.627 LAYER MTL1  ;
	END SCEN
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER MTL1 ;
			RECT 38.9 8.58 39.92 11.22 ;
			RECT 39.28 2.16 39.92 11.22 ;
			RECT 39.2 2.16 39.92 2.8 ;

		END 

		ANTENNADIFFAREA 3.828 LAYER MTL1  ;
	END Q
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 40.32 13.68 ;
			RECT 37.44 8.58 38.08 13.68 ;
			RECT 35.56 10.7 36.2 13.68 ;
			RECT 28.64 8.58 29.28 13.68 ;
			RECT 25.68 9.36 26.32 13.68 ;
			RECT 19.64 10.7 20.28 13.68 ;
			RECT 13.24 10.94 13.88 13.68 ;
			RECT 9.44 11.66 10.08 13.68 ;
			RECT 1 10.9 1.64 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 40.32 1.46 ;
			RECT 37.8 -0.48 38.44 2.76 ;
			RECT 33.48 -0.48 34.12 3.7 ;
			RECT 28.68 -0.48 29.32 3.44 ;
			RECT 25.16 -0.48 25.8 2.06 ;
			RECT 20.18 -0.48 20.82 1.78 ;
			RECT 13.16 -0.48 13.8 1.62 ;
			RECT 9.56 -0.48 10.2 2.26 ;
			RECT 1 -0.48 1.64 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1 2.78 5.04 3.26 ;
			RECT 1 2.78 1.64 3.9 ;
			RECT 4.44 2.78 5.04 5.62 ;
			RECT 4.44 3.98 5.56 5.62 ;
			RECT 4.44 7.86 6.66 8.5 ;
			RECT 4.44 2.78 4.92 10.2 ;
			RECT 1 9.54 4.92 10.2 ;
			RECT 11.72 3.14 12.36 4.42 ;
			RECT 8.72 3.78 12.36 4.42 ;
			RECT 11.2 3.78 11.68 10.14 ;
			RECT 15.24 8.4 15.88 9.42 ;
			RECT 11.2 8.94 15.88 9.42 ;
			RECT 11.2 8.94 11.72 10.14 ;
			RECT 11.08 9.5 11.72 10.14 ;
			RECT 12.24 9.94 15.24 10.42 ;
			RECT 14.76 9.94 15.24 11.22 ;
			RECT 5.48 9.4 6.12 11.14 ;
			RECT 12.24 9.94 12.72 11.14 ;
			RECT 5.48 10.66 12.72 11.14 ;
			RECT 14.76 10.58 16.44 11.22 ;
			RECT 15.8 1.98 16.44 2.62 ;
			RECT 10.72 2.14 16.44 2.62 ;
			RECT 10.72 2.14 11.2 3.26 ;
			RECT 5.56 2.78 11.2 3.26 ;
			RECT 5.56 2.78 6.2 3.46 ;
			RECT 18.18 3.3 18.82 4.94 ;
			RECT 16.84 4.46 18.82 4.94 ;
			RECT 16.84 4.46 17.32 9.04 ;
			RECT 16.68 8.4 17.32 9.04 ;
			RECT 17.52 1.98 18.2 2.78 ;
			RECT 17.52 2.3 20.82 2.78 ;
			RECT 20.2 2.3 20.82 10.04 ;
			RECT 20.2 2.94 21.28 3.58 ;
			RECT 20.2 2.94 20.84 10.04 ;
			RECT 17.2 9.56 20.84 10.04 ;
			RECT 17.2 9.56 17.84 11.22 ;
			RECT 21.8 1.98 22.46 11.22 ;
			RECT 21.08 10.56 22.46 11.22 ;
			RECT 23.64 1.98 24.28 3.06 ;
			RECT 23.16 2.58 25.84 3.06 ;
			RECT 25.36 2.58 25.84 3.78 ;
			RECT 25.36 3.14 27.16 3.78 ;
			RECT 23.16 2.58 23.64 10 ;
			RECT 23.16 6.98 23.8 10 ;
			RECT 23.16 9.36 24.92 10 ;
			RECT 26.92 1.98 28.16 2.62 ;
			RECT 27.68 1.98 28.16 6.22 ;
			RECT 27.12 5.58 28.78 6.22 ;
			RECT 27.12 5.58 27.76 10.12 ;
			RECT 30.08 2.8 30.72 11.22 ;
			RECT 34.92 8.54 36.56 9.18 ;
			RECT 34.92 8.54 35.56 10.18 ;
			RECT 34.92 1.98 36.76 2.62 ;
			RECT 34.92 1.98 35.56 6.58 ;
			RECT 36.12 3.44 38.76 4.08 ;
			RECT 36.12 3.44 36.6 8.02 ;
			RECT 31.48 7.38 38.6 8.02 ;
			RECT 31.48 2.8 32.12 11.22 ;
			RECT 31.48 10.58 33.56 11.22 ;

	END

END DFCH

MACRO DEL_50NS_RC
	CLASS CORE ;
	FOREIGN DEL_50NS_RC 0 0  ;
	ORIGIN 0 0 ;
	SIZE 46.08 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN DIN
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.605 LAYER MTL1  ;
	END DIN
	PIN DOUT
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 45.04 1.98 45.68 11.22 ;
			RECT 43.52 1.98 45.68 4.06 ;

		END 

		ANTENNADIFFAREA 5.491 LAYER MTL1  ;
	END DOUT
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 46.08 13.68 ;
			RECT 43.16 5.42 43.8 10.66 ;
			RECT 42.8 10.14 43.44 13.68 ;
			RECT 33.3 8.58 33.94 13.68 ;
			RECT 4.7 8.58 5.34 13.68 ;
			RECT 1.84 10.26 2.48 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 46.08 1.46 ;
			RECT 41.92 -0.48 42.72 3.98 ;
			RECT 41.92 -0.48 42.56 9.62 ;
			RECT 34.12 -0.48 34.76 2.54 ;
			RECT 32.48 -0.48 33.12 4.26 ;
			RECT 27.16 -0.48 27.8 4.26 ;
			RECT 1.72 -0.48 2.36 2.64 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1.68 3.66 2.7 4.3 ;
			RECT 2.06 3.66 2.7 9.74 ;
			RECT 0.4 9.26 2.7 9.74 ;
			RECT 0.4 9.26 1.04 11.22 ;
			RECT 3.2 1.98 5.86 2.62 ;
			RECT 3.2 1.98 3.92 2.64 ;
			RECT 3.28 1.98 3.92 11.22 ;
			RECT 3.22 9.28 3.92 11.22 ;
			RECT 28.04 4.78 34.16 7.98 ;
			RECT 5.58 7.34 34.16 7.98 ;
			RECT 39.04 2.96 39.68 5.7 ;
			RECT 36.64 5.06 39.68 5.7 ;
			RECT 36.64 5.06 37.28 10.22 ;
			RECT 40.68 2.96 41.32 6.7 ;
			RECT 39.4 6.22 41.32 6.7 ;
			RECT 39.4 6.22 40.04 10.22 ;
			RECT 35.64 3.34 36.84 3.98 ;
			RECT 35.64 3.34 36.12 11.22 ;
			RECT 41.4 10.14 42.04 11.22 ;
			RECT 35.64 10.74 42.04 11.22 ;

	END

END DEL_50NS_RC

MACRO DEL_30NS_RC
	CLASS CORE ;
	FOREIGN DEL_30NS_RC 0 0  ;
	ORIGIN 0 0 ;
	SIZE 46.08 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN DIN
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.605 LAYER MTL1  ;
	END DIN
	PIN DOUT
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 45.04 1.98 45.68 11.22 ;
			RECT 43.52 1.98 45.68 4.06 ;

		END 

		ANTENNADIFFAREA 5.491 LAYER MTL1  ;
	END DOUT
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 46.08 13.68 ;
			RECT 43.16 5.42 43.8 10.66 ;
			RECT 42.8 10.14 43.44 13.68 ;
			RECT 33.3 8.58 33.94 13.68 ;
			RECT 4.7 8.58 5.34 13.68 ;
			RECT 1.84 10.26 2.48 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 46.08 1.46 ;
			RECT 41.92 -0.48 42.72 3.98 ;
			RECT 41.92 -0.48 42.56 9.62 ;
			RECT 34.12 -0.48 34.76 2.54 ;
			RECT 32.48 -0.48 33.12 4.26 ;
			RECT 27.16 -0.48 27.8 4.26 ;
			RECT 1.72 -0.48 2.36 2.64 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1.68 3.66 2.7 4.3 ;
			RECT 2.06 3.66 2.7 9.74 ;
			RECT 0.4 9.26 2.7 9.74 ;
			RECT 0.4 9.26 1.04 11.22 ;
			RECT 3.2 1.98 5.86 2.62 ;
			RECT 3.2 1.98 3.92 2.64 ;
			RECT 3.28 1.98 3.92 11.22 ;
			RECT 3.22 9.28 3.92 11.22 ;
			RECT 5.22 5.9 5.86 7.98 ;
			RECT 28.04 4.78 34.16 7.98 ;
			RECT 5.22 7.34 34.16 7.98 ;
			RECT 39.04 2.96 39.68 5.7 ;
			RECT 36.64 5.06 39.68 5.7 ;
			RECT 36.64 5.06 37.28 10.22 ;
			RECT 40.68 2.96 41.32 6.7 ;
			RECT 39.4 6.22 41.32 6.7 ;
			RECT 39.4 6.22 40.04 10.22 ;
			RECT 35.64 3.34 36.84 3.98 ;
			RECT 35.64 3.34 36.12 11.22 ;
			RECT 41.4 10.14 42.04 11.22 ;
			RECT 35.64 10.74 42.04 11.22 ;

	END

END DEL_30NS_RC

MACRO DEL_20NS_RC
	CLASS CORE ;
	FOREIGN DEL_20NS_RC 0 0  ;
	ORIGIN 0 0 ;
	SIZE 33.12 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN DIN
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.605 LAYER MTL1  ;
	END DIN
	PIN DOUT
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 32.08 1.98 32.72 11.22 ;
			RECT 30.56 1.98 32.72 4.06 ;

		END 

		ANTENNADIFFAREA 5.491 LAYER MTL1  ;
	END DOUT
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 33.12 13.68 ;
			RECT 30.2 5.42 30.84 10.66 ;
			RECT 29.84 10.14 30.48 13.68 ;
			RECT 20.24 8.58 20.88 13.68 ;
			RECT 4.7 8.58 5.34 13.68 ;
			RECT 1.84 10.26 2.48 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 33.12 1.46 ;
			RECT 28.96 -0.48 29.76 3.98 ;
			RECT 28.96 -0.48 29.6 9.62 ;
			RECT 21.16 -0.48 21.8 2.54 ;
			RECT 1.72 -0.48 2.36 2.64 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1.68 3.66 2.7 4.3 ;
			RECT 2.06 3.66 2.7 9.74 ;
			RECT 0.4 9.26 2.7 9.74 ;
			RECT 0.4 9.26 1.04 11.22 ;
			RECT 3.2 1.98 5.62 2.62 ;
			RECT 3.2 1.98 3.92 2.64 ;
			RECT 3.28 1.98 3.92 11.22 ;
			RECT 3.22 9.28 3.92 11.22 ;
			RECT 4.44 5.94 5.08 7.98 ;
			RECT 21.52 3.62 22.16 7.98 ;
			RECT 4.44 7.34 22.16 7.98 ;
			RECT 26.08 2.96 26.72 5.7 ;
			RECT 23.68 5.06 26.72 5.7 ;
			RECT 23.68 5.06 24.32 10.22 ;
			RECT 27.72 2.96 28.36 6.7 ;
			RECT 26.44 6.22 28.36 6.7 ;
			RECT 26.44 6.22 27.08 10.22 ;
			RECT 22.68 3.34 23.88 3.98 ;
			RECT 22.68 3.34 23.16 11.22 ;
			RECT 28.44 10.14 29.08 11.22 ;
			RECT 22.68 10.74 29.08 11.22 ;

	END

END DEL_20NS_RC

MACRO DEL_10NS_RC
	CLASS CORE ;
	FOREIGN DEL_10NS_RC 0 0  ;
	ORIGIN 0 0 ;
	SIZE 33.12 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN DIN
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.605 LAYER MTL1  ;
	END DIN
	PIN DOUT
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 32.08 1.98 32.72 11.22 ;
			RECT 30.56 1.98 32.72 4.06 ;

		END 

		ANTENNADIFFAREA 5.491 LAYER MTL1  ;
	END DOUT
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 33.12 13.68 ;
			RECT 30.2 5.42 30.84 10.66 ;
			RECT 29.84 10.14 30.48 13.68 ;
			RECT 20.24 8.58 20.88 13.68 ;
			RECT 4.7 8.58 5.34 13.68 ;
			RECT 1.84 10.26 2.48 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 33.12 1.46 ;
			RECT 28.96 -0.48 29.76 3.98 ;
			RECT 28.96 -0.48 29.6 9.62 ;
			RECT 21.16 -0.48 21.8 2.54 ;
			RECT 1.72 -0.48 2.36 2.64 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1.68 3.66 2.7 4.3 ;
			RECT 2.06 3.66 2.7 9.74 ;
			RECT 0.4 9.26 2.7 9.74 ;
			RECT 0.4 9.26 1.04 11.22 ;
			RECT 3.2 1.98 5.76 2.62 ;
			RECT 3.2 1.98 3.92 2.64 ;
			RECT 3.28 1.98 3.92 11.22 ;
			RECT 3.22 9.28 3.92 11.22 ;
			RECT 5.12 5.9 5.76 7.98 ;
			RECT 20.56 3.96 21.2 7.98 ;
			RECT 5.12 7.34 21.2 7.98 ;
			RECT 26.08 2.96 26.72 5.7 ;
			RECT 23.68 5.06 26.72 5.7 ;
			RECT 23.68 5.06 24.32 10.22 ;
			RECT 27.72 2.96 28.36 6.7 ;
			RECT 26.44 6.22 28.36 6.7 ;
			RECT 26.44 6.22 27.08 10.22 ;
			RECT 22.68 3.34 23.88 3.98 ;
			RECT 22.68 3.34 23.16 11.22 ;
			RECT 28.44 10.14 29.08 11.22 ;
			RECT 22.68 10.74 29.08 11.22 ;

	END

END DEL_10NS_RC

MACRO DEL3RC
	CLASS CORE ;
	FOREIGN DEL3RC 0 0  ;
	ORIGIN 0 0 ;
	SIZE 17.28 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.749 LAYER MTL1  ;
	END A
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 16.24 1.98 16.88 11.22 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 17.28 13.68 ;
			RECT 14.76 10.22 15.4 13.68 ;
			RECT 1.8 10.7 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 17.28 1.46 ;
			RECT 14.8 -0.48 15.44 2.62 ;
			RECT 0.88 -0.48 1.52 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1 3.26 2.76 3.9 ;
			RECT 2.28 5.62 3.92 6.26 ;
			RECT 2.28 3.26 2.76 10.18 ;
			RECT 0.4 9.7 2.76 10.18 ;
			RECT 0.4 9.7 1.04 11.22 ;

	END

END DEL3RC

MACRO DEL20
	CLASS CORE ;
	FOREIGN DEL20 0 0  ;
	ORIGIN 0 0 ;
	SIZE 33.12 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 4.96 1.04 6.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.648 LAYER MTL1  ;
	END A
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 32.08 2 32.72 10.88 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 33.12 13.68 ;
			RECT 30.68 10.3 31.32 13.68 ;
			RECT 21.48 10.7 22.12 13.68 ;
			RECT 11.64 10.7 12.28 13.68 ;
			RECT 1.8 10.7 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 33.12 1.46 ;
			RECT 30.68 -0.48 31.32 2.64 ;
			RECT 22.64 -0.48 23.28 2.5 ;
			RECT 12.38 -0.48 13.02 2.5 ;
			RECT 2.04 -0.48 2.7 2.5 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 1.98 1.04 3.5 ;
			RECT 0.4 3.02 3.92 3.5 ;
			RECT 3.28 3.02 3.92 10.18 ;
			RECT 0.4 9.7 3.92 10.18 ;
			RECT 0.4 9.7 1.04 11.22 ;
			RECT 6.5 1.98 7.14 4.1 ;
			RECT 6.16 3.46 8.32 4.1 ;
			RECT 6.16 3.46 6.64 11.22 ;
			RECT 6 10.58 6.64 11.22 ;
			RECT 7.9 1.98 9.6 2.62 ;
			RECT 9.12 3.46 13.62 4.1 ;
			RECT 9.12 1.98 9.6 5.1 ;
			RECT 7.44 4.62 9.6 5.1 ;
			RECT 7.44 4.62 7.92 11.22 ;
			RECT 7.44 10.58 8.08 11.22 ;
			RECT 16.82 1.98 17.68 2.62 ;
			RECT 17.04 1.98 17.68 4.98 ;
			RECT 17.04 4.34 18.68 4.98 ;
			RECT 18.2 4.34 18.68 10.06 ;
			RECT 15.84 9.58 18.68 10.06 ;
			RECT 15.84 9.58 16.48 11.22 ;
			RECT 18.4 3.18 23.92 3.82 ;
			RECT 19.2 3.18 23.92 4.1 ;
			RECT 19.2 3.18 19.68 11.22 ;
			RECT 17.28 10.58 19.68 11.22 ;
			RECT 26.36 3.18 28.56 4.82 ;
			RECT 26.36 3.18 26.9 11.22 ;
			RECT 25.68 10.58 26.9 11.22 ;
			RECT 28.32 2 29.8 2.64 ;
			RECT 29.32 3.22 31.56 4.86 ;
			RECT 29.32 2 29.8 11.22 ;
			RECT 28.32 10.58 29.8 11.22 ;

	END

END DEL20

MACRO DEL10
	CLASS CORE ;
	FOREIGN DEL10 0 0  ;
	ORIGIN 0 0 ;
	SIZE 27.36 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 4.96 1.04 6.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.648 LAYER MTL1  ;
	END A
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 26.32 2 26.96 10.88 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 27.36 13.68 ;
			RECT 24.92 10.3 25.56 13.68 ;
			RECT 16.84 10.7 17.48 13.68 ;
			RECT 9.32 10.7 9.96 13.68 ;
			RECT 1.8 10.7 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 27.36 1.46 ;
			RECT 24.92 -0.48 25.56 2.64 ;
			RECT 18.04 -0.48 18.68 2.5 ;
			RECT 10.06 -0.48 10.7 2.5 ;
			RECT 2.04 -0.48 2.7 2.5 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 1.98 1.04 3.5 ;
			RECT 0.4 3.02 3.92 3.5 ;
			RECT 3.28 3.02 3.92 10.18 ;
			RECT 0.4 9.7 3.92 10.18 ;
			RECT 0.4 9.7 1.04 11.22 ;
			RECT 5.34 1.98 5.98 4.1 ;
			RECT 4.8 3.46 7.16 4.1 ;
			RECT 4.8 3.46 5.28 11.22 ;
			RECT 4.8 10.58 5.48 11.22 ;
			RECT 6.74 1.98 8.16 2.62 ;
			RECT 7.68 3.46 11.3 4.1 ;
			RECT 7.68 1.98 8.16 5.1 ;
			RECT 6.44 4.62 8.16 5.1 ;
			RECT 6.44 4.62 6.92 11.22 ;
			RECT 6.28 10.58 6.92 11.22 ;
			RECT 13.34 1.98 14.32 2.62 ;
			RECT 13.68 1.98 14.32 4.98 ;
			RECT 13.68 4.34 15.32 4.98 ;
			RECT 14.68 4.34 15.32 10.06 ;
			RECT 12.36 9.58 15.32 10.06 ;
			RECT 12.36 9.58 13 11.22 ;
			RECT 14.96 3.18 19.28 3.82 ;
			RECT 15.84 3.18 19.28 4.1 ;
			RECT 15.84 3.18 16.32 11.22 ;
			RECT 13.8 10.58 16.32 11.22 ;
			RECT 21.12 3.18 22.76 4.82 ;
			RECT 21.12 3.18 21.76 11.22 ;
			RECT 19.88 10.58 21.76 11.22 ;
			RECT 22.56 2 24 2.64 ;
			RECT 23.52 3.22 25.8 4.86 ;
			RECT 23.52 2 24 11.22 ;
			RECT 22.56 10.58 24 11.22 ;

	END

END DEL10

MACRO DECAP8
	CLASS CORE SPACER ;
	FOREIGN DECAP8 0 0  ;
	ORIGIN 0 0 ;
	SIZE 11.52 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 11.52 13.68 ;
			RECT 0.72 10.7 10.8 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 11.52 1.46 ;
			RECT 3.28 -0.48 8.24 1.82 ;

		END 

	END gndd!

END DECAP8

MACRO DECAP4
	CLASS CORE SPACER ;
	FOREIGN DECAP4 0 0  ;
	ORIGIN 0 0 ;
	SIZE 5.76 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 5.76 13.68 ;
			RECT 1.06 10.7 4.7 13.68 ;
			RECT 1.06 8.22 4.7 8.86 ;
			RECT 2.54 8.22 3.22 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 5.76 1.46 ;
			RECT 0.32 -0.48 5.44 1.82 ;

		END 

	END gndd!

END DECAP4

MACRO DECAP16
	CLASS CORE SPACER ;
	FOREIGN DECAP16 0 0  ;
	ORIGIN 0 0 ;
	SIZE 23.04 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 23.04 13.68 ;
			RECT 0.72 10.7 22.32 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 23.04 1.46 ;
			RECT 3.26 -0.48 19.74 1.82 ;

		END 

	END gndd!

END DECAP16

MACRO BF8
	CLASS CORE ;
	FOREIGN BF8 0 0  ;
	ORIGIN 0 0 ;
	SIZE 27.36 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.96 3.48 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 5.76 LAYER MTL1  ;
	END A
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 23.88 2.82 26.82 8.04 ;
			RECT 24.76 1.98 25.4 11.22 ;
			RECT 7.88 6.82 25.4 8.06 ;
			RECT 7.96 2.8 25.4 3.72 ;
			RECT 21.96 6.82 22.6 11.22 ;
			RECT 21.96 1.98 22.6 3.72 ;
			RECT 19.12 6.82 19.84 11.22 ;
			RECT 19.16 1.98 19.8 3.72 ;
			RECT 16.36 1.98 17 3.72 ;
			RECT 16.32 6.82 16.96 11.22 ;
			RECT 13.56 1.98 14.2 3.72 ;
			RECT 13.52 6.82 14.16 11.22 ;
			RECT 10.68 6.82 11.4 11.22 ;
			RECT 7.96 2.78 11.4 3.72 ;
			RECT 10.76 1.98 11.4 3.72 ;
			RECT 7.88 6.82 8.6 11.22 ;
			RECT 7.96 1.98 8.6 3.72 ;

		END 

		ANTENNADIFFAREA 32.614 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 27.36 13.68 ;
			RECT 26.16 8.56 26.8 13.68 ;
			RECT 23.36 8.58 24 13.68 ;
			RECT 20.52 8.58 21.24 13.68 ;
			RECT 17.68 8.58 18.4 13.68 ;
			RECT 14.92 8.58 15.56 13.68 ;
			RECT 12.12 8.58 12.76 13.68 ;
			RECT 9.3 8.58 9.96 13.68 ;
			RECT 6.44 8.58 7.08 13.68 ;
			RECT 3.64 8.44 4.28 13.68 ;
			RECT 0.84 8.44 1.48 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 27.36 1.46 ;
			RECT 26.16 -0.48 26.8 2.28 ;
			RECT 23.36 -0.48 24 2.28 ;
			RECT 20.56 -0.48 21.2 2.28 ;
			RECT 17.76 -0.48 18.4 2.28 ;
			RECT 14.96 -0.48 15.6 2.28 ;
			RECT 12.16 -0.48 12.8 2.28 ;
			RECT 9.36 -0.48 10 2.26 ;
			RECT 6.56 -0.48 7.2 2.54 ;
			RECT 3.64 -0.48 4.28 2.54 ;
			RECT 0.84 -0.48 1.48 2.62 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 2.24 1.98 2.88 3.86 ;
			RECT 2.24 3.06 5.68 3.86 ;
			RECT 4.76 3.06 5.68 7.92 ;
			RECT 4.76 4.48 21.62 5.84 ;
			RECT 4.76 4.48 6.08 7.92 ;
			RECT 2.24 7.14 6.08 7.92 ;
			RECT 2.24 7.14 2.88 11.22 ;
			RECT 5.04 1.98 5.68 11.22 ;

	END

END BF8

MACRO BF5
	CLASS CORE ;
	FOREIGN BF5 0 0  ;
	ORIGIN 0 0 ;
	SIZE 12.96 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 3.211 LAYER MTL1  ;
	END A
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 10.28 7.58 10.92 11.22 ;
			RECT 4.64 7.58 10.92 8.06 ;
			RECT 7.44 7.58 8.16 11.22 ;
			RECT 3.28 3.64 6.72 4.28 ;
			RECT 6.08 1.98 6.72 4.28 ;
			RECT 4.64 7.58 5.36 11.22 ;
			RECT 4.72 3.64 5.36 11.22 ;
			RECT 3.28 1.98 3.92 4.28 ;

		END 

		ANTENNADIFFAREA 15.027 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 12.96 13.68 ;
			RECT 11.8 8.58 12.44 13.68 ;
			RECT 8.88 8.58 9.52 13.68 ;
			RECT 6.06 8.58 6.72 13.68 ;
			RECT 3.2 8.58 3.84 13.68 ;
			RECT 0.4 8.44 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 12.96 1.46 ;
			RECT 7.48 -0.48 8.12 3.78 ;
			RECT 4.68 -0.48 5.32 3.1 ;
			RECT 1.8 -0.48 2.44 3.58 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 1.98 1.04 4.76 ;
			RECT 0.4 4.28 2.76 4.76 ;
			RECT 2.28 4.28 2.76 5.44 ;
			RECT 2.28 4.8 4.2 5.44 ;
			RECT 2.72 4.8 3.2 8.06 ;
			RECT 1.8 7.54 3.2 8.06 ;
			RECT 1.8 7.54 2.44 11.22 ;

	END

END BF5

MACRO BF4
	CLASS CORE ;
	FOREIGN BF4 0 0  ;
	ORIGIN 0 0 ;
	SIZE 10.08 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.462 LAYER MTL1  ;
	END A
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.52 7.76 8.16 11.22 ;
			RECT 3.28 7.76 8.16 8.24 ;
			RECT 4.62 9.54 5.36 11.22 ;
			RECT 4.72 6.28 5.36 11.22 ;
			RECT 3.28 7.6 5.36 8.24 ;
			RECT 3.44 6.28 5.36 8.24 ;
			RECT 3.44 1.98 3.92 8.24 ;
			RECT 3.28 1.98 3.92 4.3 ;

		END 

		ANTENNADIFFAREA 10.138 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 10.08 13.68 ;
			RECT 8.92 9.36 9.56 13.68 ;
			RECT 6.04 9.7 6.7 13.68 ;
			RECT 3.2 9.58 3.84 13.68 ;
			RECT 0.4 9.58 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 10.08 1.46 ;
			RECT 4.68 -0.48 5.32 4.42 ;
			RECT 1.8 -0.48 2.44 3.58 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 2.28 1.04 4.76 ;
			RECT 0.4 4.28 2.76 4.76 ;
			RECT 2.2 4.28 2.76 6.54 ;
			RECT 2.2 4.9 2.92 6.54 ;
			RECT 2.2 4.28 2.68 11.22 ;
			RECT 1.8 9.58 2.68 11.22 ;

	END

END BF4

MACRO BF3
	CLASS CORE ;
	FOREIGN BF3 0 0  ;
	ORIGIN 0 0 ;
	SIZE 8.64 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 5.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.901 LAYER MTL1  ;
	END A
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.52 7.44 8.16 11.22 ;
			RECT 4.72 7.44 8.16 8.08 ;
			RECT 3.68 3.14 6.72 3.62 ;
			RECT 6.08 1.98 6.72 3.62 ;
			RECT 4.72 3.14 5.36 8.24 ;
			RECT 4.62 7.74 5.34 11.22 ;
			RECT 3.68 1.98 4.16 3.62 ;
			RECT 3.28 1.98 4.16 2.64 ;

		END 

		ANTENNADIFFAREA 8.73 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 8.64 13.68 ;
			RECT 6.04 8.6 6.7 13.68 ;
			RECT 3.2 9.58 3.84 13.68 ;
			RECT 0.4 9.58 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 8.64 1.46 ;
			RECT 7.48 -0.48 8.12 2.62 ;
			RECT 4.68 -0.48 5.32 2.62 ;
			RECT 1.8 -0.48 2.44 2.64 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 2.28 1.04 3.64 ;
			RECT 0.4 3.16 3.16 3.64 ;
			RECT 2.68 3.16 3.16 4.62 ;
			RECT 2.68 4.14 4.2 4.62 ;
			RECT 3.56 4.14 4.2 5.92 ;
			RECT 3.56 4.14 4.04 9.06 ;
			RECT 1.8 8.58 4.04 9.06 ;
			RECT 1.8 8.58 2.44 11.22 ;

	END

END BF3

MACRO BF2
	CLASS CORE ;
	FOREIGN BF2 0 0  ;
	ORIGIN 0 0 ;
	SIZE 5.76 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.138 LAYER MTL1  ;
	END A
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.24 9.52 3.92 11.22 ;
			RECT 3.28 1.98 3.92 11.22 ;

		END 

		ANTENNADIFFAREA 4.557 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 5.76 13.68 ;
			RECT 4.64 9.44 5.3 13.68 ;
			RECT 1.8 9.44 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 5.76 1.46 ;
			RECT 1.8 -0.48 2.44 2.86 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 1.98 1.04 3.86 ;
			RECT 0.4 3.38 2.76 3.86 ;
			RECT 2.12 3.38 2.76 8.92 ;
			RECT 0.4 8.44 2.76 8.92 ;
			RECT 0.4 8.44 1.04 11.22 ;

	END

END BF2

MACRO BF
	CLASS CORE ;
	FOREIGN BF 0 0  ;
	ORIGIN 0 0 ;
	SIZE 4.32 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 5.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.605 LAYER MTL1  ;
	END A
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.22 9.28 3.92 11.22 ;
			RECT 3.28 1.98 3.92 11.22 ;
			RECT 3.2 1.98 3.92 2.64 ;

		END 

		ANTENNADIFFAREA 3.168 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 4.32 13.68 ;
			RECT 1.84 10.26 2.48 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 4.32 1.46 ;
			RECT 1.72 -0.48 2.36 2.64 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1.68 3.66 2.7 4.3 ;
			RECT 2.06 3.66 2.7 9.74 ;
			RECT 0.4 9.26 2.7 9.74 ;
			RECT 0.4 9.26 1.04 11.22 ;

	END

END BF

MACRO ANTENNA
	CLASS CORE ANTENNACELL ;
	FOREIGN ANTENNA 0 0  ;
	ORIGIN 0 0 ;
	SIZE 1.44 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 2.32 1.04 2.96 ;

		END 

		ANTENNADIFFAREA 0.518 LAYER MTL1  ;
	END A
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 1.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 1.44 1.46 ;

		END 

	END gndd!

END ANTENNA

MACRO AND4XL
	CLASS CORE ;
	FOREIGN AND4XL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 8.64 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 8.92 1.04 9.56 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.619 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 7.6 2.48 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.619 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.28 3.92 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.619 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 3.96 5.36 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.619 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.48 9.02 8.24 11.22 ;
			RECT 7.6 1.98 8.24 11.22 ;
			RECT 7 1.98 8.24 2.62 ;

		END 

		ANTENNADIFFAREA 1.672 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 8.64 13.68 ;
			RECT 6.04 10.7 6.68 13.68 ;
			RECT 3.24 10.7 3.88 13.68 ;
			RECT 0.44 10.7 1.08 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 8.64 1.46 ;
			RECT 5.36 -0.48 6 2.44 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.84 1.98 1.48 3.44 ;
			RECT 0.84 2.96 6.48 3.44 ;
			RECT 6 3.14 7.08 3.8 ;
			RECT 6.44 3.14 7.08 4.8 ;
			RECT 6.44 3.14 6.92 10.18 ;
			RECT 1.84 9.7 6.92 10.18 ;
			RECT 1.84 9.7 2.48 11.22 ;
			RECT 4.64 9.7 5.28 11.22 ;

	END

END AND4XL

MACRO AND4
	CLASS CORE ;
	FOREIGN AND4 0 0  ;
	ORIGIN 0 0 ;
	SIZE 8.64 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 8.92 1.04 9.56 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.821 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 7.6 2.48 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.821 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.28 3.92 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.821 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 3.96 5.36 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.821 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.48 9.02 8.24 11.22 ;
			RECT 7.6 1.98 8.24 11.22 ;
			RECT 6.88 1.98 8.24 2.62 ;

		END 

		ANTENNADIFFAREA 3.322 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 8.64 13.68 ;
			RECT 6.04 10.7 6.68 13.68 ;
			RECT 3.24 10.7 3.88 13.68 ;
			RECT 0.44 10.7 1.08 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 8.64 1.46 ;
			RECT 5.24 -0.48 5.88 2.38 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.84 1.98 4.72 2.46 ;
			RECT 0.84 1.98 1.48 2.62 ;
			RECT 4.24 1.98 4.72 3.38 ;
			RECT 4.24 2.9 6.36 3.38 ;
			RECT 5.88 3.14 7.08 3.62 ;
			RECT 6.44 3.14 7.08 4.8 ;
			RECT 6.44 3.14 6.92 10.18 ;
			RECT 1.84 9.7 6.92 10.18 ;
			RECT 1.84 9.7 2.48 11.22 ;
			RECT 4.64 9.7 5.28 11.22 ;

	END

END AND4

MACRO AND3XL
	CLASS CORE ;
	FOREIGN AND3XL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 7.54 1.04 9.18 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.562 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 3.98 2.48 5.62 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.562 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.28 3.92 7.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.562 LAYER MTL1  ;
	END C
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.04 10.24 6.8 11.22 ;
			RECT 6.16 1.98 6.8 11.22 ;
			RECT 5.68 1.98 6.8 2.62 ;

		END 

		ANTENNADIFFAREA 1.614 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 4.6 10.7 5.24 13.68 ;
			RECT 1.8 10.7 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 4.04 -0.48 4.68 2.62 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 1.98 1.04 3.44 ;
			RECT 0.4 2.96 3.52 3.44 ;
			RECT 3.04 3.14 5.64 3.62 ;
			RECT 5 3.14 5.64 4.8 ;
			RECT 5 3.14 5.48 10.18 ;
			RECT 0.4 9.7 5.48 10.18 ;
			RECT 0.4 9.7 1.04 11.22 ;
			RECT 3.2 9.7 3.84 11.22 ;

	END

END AND3XL

MACRO AND32OXL
	CLASS CORE ;
	FOREIGN AND32OXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 8.64 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 7.6 1.04 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.037 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.037 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 3.96 3.92 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.037 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 3.96 6.8 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.965 LAYER MTL1  ;
	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 6.28 5.36 7.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.965 LAYER MTL1  ;
	END E
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6 9.42 8.24 10.06 ;
			RECT 7.6 1.98 8.24 10.06 ;
			RECT 0.4 2.96 8.24 3.44 ;
			RECT 6.44 1.98 8.24 3.44 ;
			RECT 0.4 1.98 1.04 3.44 ;

		END 

		ANTENNADIFFAREA 3.698 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 8.64 13.68 ;
			RECT 3.2 9.46 3.84 13.68 ;
			RECT 0.4 9.42 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 8.64 1.46 ;
			RECT 3.8 -0.48 4.44 2.44 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1.8 8.46 5.24 8.94 ;
			RECT 4.6 8.46 5.24 11.22 ;
			RECT 1.8 8.46 2.44 11.18 ;
			RECT 4.6 10.58 8.04 11.22 ;

	END

END AND32OXL

MACRO AND32O
	CLASS CORE ;
	FOREIGN AND32O 0 0  ;
	ORIGIN 0 0 ;
	SIZE 12.96 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.84 4.96 2.48 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.376 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.22 3.92 7.86 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.376 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 6.22 6.8 7.86 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.376 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 10.48 5.28 11.12 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.261 LAYER MTL1  ;
	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 4.96 8.24 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.261 LAYER MTL1  ;
	END E
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.72 10.58 12.56 11.22 ;
			RECT 11.92 1.98 12.56 11.22 ;
			RECT 6.32 1.98 12.56 2.62 ;
			RECT 4.16 2.9 6.8 3.38 ;
			RECT 6.32 1.98 6.8 3.38 ;
			RECT 4.16 1.98 4.64 3.38 ;
			RECT 1.76 1.98 4.64 2.62 ;

		END 

		ANTENNADIFFAREA 8.086 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 12.96 13.68 ;
			RECT 4.92 9.7 5.56 13.68 ;
			RECT 0.8 10.58 2.76 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 12.96 1.46 ;
			RECT 5.16 -0.48 5.8 2.38 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 2.12 8.7 10.76 9.18 ;
			RECT 2.12 8.7 4.4 9.82 ;
			RECT 6.08 8.7 10.76 9.82 ;
			RECT 3.52 8.7 4.4 10.82 ;
			RECT 6.08 8.7 6.96 10.82 ;

	END

END AND32O

MACRO AND31OXL
	CLASS CORE ;
	FOREIGN AND31OXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 7.6 1.04 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.037 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.037 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 3.96 3.92 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.037 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 6.28 5.36 7.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.893 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6 9.46 6.8 11.22 ;
			RECT 6.16 1.98 6.8 11.22 ;
			RECT 0.4 2.96 6.8 3.44 ;
			RECT 5.44 1.98 6.8 3.44 ;
			RECT 0.4 1.98 1.04 3.44 ;

		END 

		ANTENNADIFFAREA 3.328 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 3.2 10.08 3.84 13.68 ;
			RECT 0.4 9.46 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 3.8 -0.48 4.44 2.44 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1.8 8.76 5.24 9.24 ;
			RECT 1.8 8.76 2.44 11.22 ;
			RECT 4.6 8.76 5.24 11.22 ;

	END

END AND31OXL

MACRO AND31O
	CLASS CORE ;
	FOREIGN AND31O 0 0  ;
	ORIGIN 0 0 ;
	SIZE 10.08 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.02 2.48 5.66 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.376 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.22 3.92 7.86 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.376 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 6.22 6.8 7.86 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.376 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 3.96 8.24 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.059 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.72 10.58 9.68 11.22 ;
			RECT 9.04 1.98 9.68 11.22 ;
			RECT 6.6 1.98 9.68 2.62 ;
			RECT 1.76 2.9 7.24 3.38 ;
			RECT 6.6 1.98 7.24 3.38 ;
			RECT 1.76 1.98 2.4 3.38 ;

		END 

		ANTENNADIFFAREA 6.706 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 10.08 13.68 ;
			RECT 4.92 9.7 5.56 13.68 ;
			RECT 0.8 10.58 2.76 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 10.08 1.46 ;
			RECT 5.16 -0.48 5.8 2.38 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 2.12 8.7 8.36 9.18 ;
			RECT 2.12 8.7 4.4 9.82 ;
			RECT 6.08 8.7 8.36 9.82 ;
			RECT 3.52 8.7 4.4 10.82 ;
			RECT 6.08 8.7 6.96 10.82 ;

	END

END AND31O

MACRO AND3
	CLASS CORE ;
	FOREIGN AND3 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 7.54 1.04 9.18 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.778 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.778 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 3.96 3.92 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.778 LAYER MTL1  ;
	END C
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.04 9.02 6.8 11.22 ;
			RECT 6.16 1.98 6.8 11.22 ;
			RECT 5.44 1.98 6.8 2.62 ;

		END 

		ANTENNADIFFAREA 3.322 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 4.6 10.7 5.24 13.68 ;
			RECT 1.8 10.7 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 3.8 -0.48 4.44 2.38 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 1.98 1.04 3.44 ;
			RECT 0.4 2.96 4.92 3.44 ;
			RECT 4.44 3.14 5.64 3.62 ;
			RECT 5 3.14 5.64 4.8 ;
			RECT 5 3.14 5.48 10.18 ;
			RECT 0.4 9.7 5.48 10.18 ;
			RECT 0.4 9.7 1.04 11.22 ;
			RECT 3.2 9.7 3.84 11.22 ;

	END

END AND3

MACRO AND2XL
	CLASS CORE ;
	FOREIGN AND2XL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 5.76 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 7.6 1.04 9.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.518 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 5.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.518 LAYER MTL1  ;
	END B
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.64 10.58 5.36 11.22 ;
			RECT 4.72 1.98 5.36 11.22 ;
			RECT 4.68 1.98 5.36 2.62 ;

		END 

		ANTENNADIFFAREA 1.614 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 5.76 13.68 ;
			RECT 3.2 10.7 3.84 13.68 ;
			RECT 0.4 10.7 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 5.76 1.46 ;
			RECT 3.04 -0.48 3.68 2.62 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 1.98 1.04 3.62 ;
			RECT 0.4 3.14 4.2 3.62 ;
			RECT 3.56 3.14 4.2 4.78 ;
			RECT 3.72 3.14 4.2 10.06 ;
			RECT 1.8 9.58 4.2 10.06 ;
			RECT 1.8 9.58 2.44 11.22 ;

	END

END AND2XL

MACRO AND2N2OXL
	CLASS CORE ;
	FOREIGN AND2N2OXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 10.08 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 3.98 2.48 5.62 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.138 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 6.6 1.04 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.138 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 6.28 6.8 7.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.21 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.34 4.96 5.36 5.62 ;
			RECT 4.34 3.98 4.98 5.62 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.21 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 8.44 9.58 9.68 11.22 ;
			RECT 9.04 3.14 9.68 11.22 ;
			RECT 6.22 3.14 9.68 3.62 ;
			RECT 6.22 1.98 6.86 3.62 ;

		END 

		ANTENNADIFFAREA 3.102 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 10.08 13.68 ;
			RECT 5.64 10.7 6.28 13.68 ;
			RECT 0.4 9.58 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 10.08 1.46 ;
			RECT 7.86 -0.48 8.5 2.62 ;
			RECT 3.68 -0.48 4.32 2.42 ;
			RECT 0.4 -0.48 1.04 2.62 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 4.24 9.7 7.68 10.18 ;
			RECT 4.24 9.7 4.92 10.78 ;
			RECT 7.04 9.7 7.68 10.78 ;
			RECT 2.04 1.98 2.68 3.44 ;
			RECT 2.04 2.94 3.48 3.44 ;
			RECT 7.4 7.76 8.18 8.42 ;
			RECT 3 2.94 3.48 9.18 ;
			RECT 7.4 7.76 7.9 9.18 ;
			RECT 2.8 8.7 7.9 9.18 ;
			RECT 2.8 8.7 3.44 10.42 ;

	END

END AND2N2OXL

MACRO AND2N2O
	CLASS CORE ;
	FOREIGN AND2N2O 0 0  ;
	ORIGIN 0 0 ;
	SIZE 11.52 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 3.96 3.92 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.138 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 7.6 1.04 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.138 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 6.28 5.36 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.462 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 4.96 8.24 6.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.462 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 10.48 1.98 11.12 11.22 ;
			RECT 8.08 2.92 11.12 3.4 ;
			RECT 8.08 1.98 8.56 3.4 ;
			RECT 6.34 1.98 8.56 2.62 ;

		END 

		ANTENNADIFFAREA 7.43 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 11.52 13.68 ;
			RECT 6.9 11.04 7.54 13.68 ;
			RECT 0.4 9.76 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 11.52 1.46 ;
			RECT 9.08 -0.48 9.72 2.4 ;
			RECT 3.68 -0.48 4.32 2.42 ;
			RECT 0.4 -0.48 1.04 2.62 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 4.16 10.04 8.94 10.52 ;
			RECT 4.16 10.04 4.84 11.16 ;
			RECT 8.3 10.04 8.94 11.22 ;
			RECT 2.04 1.98 2.68 3.42 ;
			RECT 2.04 2.94 5.64 3.42 ;
			RECT 5.14 3.14 7.56 3.64 ;
			RECT 7.08 3.14 7.56 4.42 ;
			RECT 7.08 3.92 9.8 4.42 ;
			RECT 9.32 6.18 9.96 7.84 ;
			RECT 9.32 3.92 9.8 9.52 ;
			RECT 2.8 9.04 9.8 9.52 ;
			RECT 2.8 9.04 3.44 9.68 ;

	END

END AND2N2O

MACRO AND2N1OXL
	CLASS CORE ;
	FOREIGN AND2N1OXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 7.6 1.04 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.138 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 5.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.138 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 7.6 3.92 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.138 LAYER MTL1  ;
	END C
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 5.48 8.94 6.8 11.22 ;
			RECT 6.16 3.22 6.8 11.22 ;
			RECT 4.4 3.22 6.8 3.7 ;
			RECT 4.4 3.06 5.04 3.7 ;

		END 

		ANTENNADIFFAREA 4.194 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 2.8 10 3.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 2.8 -0.48 3.44 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1.28 3.06 1.92 3.7 ;
			RECT 1.44 3.06 1.92 4.74 ;
			RECT 1.44 4.24 4.92 4.74 ;
			RECT 4.44 6.78 5.36 8.42 ;
			RECT 4.44 4.24 4.92 9.26 ;
			RECT 0.4 8.76 4.92 9.26 ;
			RECT 0.4 8.76 1.04 11.22 ;

	END

END AND2N1OXL

MACRO AND2N1O
	CLASS CORE ;
	FOREIGN AND2N1O 0 0  ;
	ORIGIN 0 0 ;
	SIZE 8.64 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 7.6 1.04 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.138 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.22 3.92 7.86 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.138 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 4.96 5.36 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.304 LAYER MTL1  ;
	END C
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 5.66 10.58 8.24 11.22 ;
			RECT 7.6 2.82 8.24 11.22 ;
			RECT 6.28 2.82 8.24 3.3 ;
			RECT 6.28 1.98 6.76 3.3 ;
			RECT 5.76 1.98 6.76 2.64 ;

		END 

		ANTENNADIFFAREA 5.844 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 8.64 13.68 ;
			RECT 2.8 10.7 3.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 8.64 1.46 ;
			RECT 7.28 -0.48 7.92 2.3 ;
			RECT 4.36 -0.48 5 2.62 ;
			RECT 1.08 -0.48 1.72 2.64 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 2.72 1.98 3.36 2.62 ;
			RECT 2.86 1.98 3.36 3.64 ;
			RECT 2.86 3.16 5.76 3.64 ;
			RECT 5.28 3.16 5.76 4.3 ;
			RECT 5.28 3.82 7.08 4.3 ;
			RECT 6.44 3.82 7.08 5.46 ;
			RECT 6.58 3.82 7.08 10.06 ;
			RECT 0.4 9.56 7.08 10.06 ;
			RECT 0.4 9.56 1.04 11.22 ;

	END

END AND2N1O

MACRO AND22OXL
	CLASS CORE ;
	FOREIGN AND22OXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 7.6 1.04 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.965 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.965 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 6.28 5.36 7.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.965 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 3.96 3.92 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.965 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.6 8.76 6.8 9.24 ;
			RECT 6.16 2.78 6.8 9.24 ;
			RECT 1.92 2.78 6.8 3.26 ;
			RECT 5.48 1.98 6.12 3.26 ;
			RECT 4.6 8.76 5.24 10.22 ;
			RECT 1.92 2.14 2.4 3.26 ;
			RECT 0.4 2.14 2.4 2.62 ;
			RECT 0.4 1.98 1.04 2.62 ;

		END 

		ANTENNADIFFAREA 3.306 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 1.8 10.02 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 2.92 -0.48 3.56 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 8.76 3.84 9.24 ;
			RECT 3.2 8.76 3.84 11.22 ;
			RECT 0.4 8.76 1.04 11.22 ;
			RECT 6 10.02 6.64 11.22 ;
			RECT 3.2 10.74 6.64 11.22 ;

	END

END AND22OXL

MACRO AND22O
	CLASS CORE ;
	FOREIGN AND22O 0 0  ;
	ORIGIN 0 0 ;
	SIZE 10.08 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 3.96 1.04 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.261 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 2.28 6.28 3.92 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.261 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 6.22 6.8 7.86 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.261 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 4.96 5.36 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.261 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 1.98 8.24 9.56 ;
			RECT 6.04 9.18 8.22 9.82 ;
			RECT 4.08 1.98 8.24 2.62 ;
			RECT 0.4 2.8 4.56 3.28 ;
			RECT 4.08 1.98 4.56 3.28 ;
			RECT 0.4 1.98 1.04 3.28 ;

		END 

		ANTENNADIFFAREA 7.589 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 10.08 13.68 ;
			RECT 3.12 10.7 3.76 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 10.08 1.46 ;
			RECT 2.92 -0.48 3.56 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1.7 9.68 5.08 10.18 ;
			RECT 4.56 9.68 5.08 11.22 ;
			RECT 1.7 9.68 2.34 11.22 ;
			RECT 0.4 10.58 2.34 11.22 ;
			RECT 4.56 10.58 8.2 11.22 ;

	END

END AND22O

MACRO AND222OXL
	CLASS CORE ;
	FOREIGN AND222OXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 10.08 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.96 2.48 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.253 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.28 3.92 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.253 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 6.28 1.04 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.253 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 4.96 5.36 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.253 LAYER MTL1  ;
	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 9.04 6.62 9.68 8.26 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.253 LAYER MTL1  ;
	END E
	PIN F
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 6.28 6.8 6.94 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.253 LAYER MTL1  ;
	END F
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.82 2.78 9.22 3.26 ;
			RECT 8.58 2.02 9.22 3.26 ;
			RECT 7.4 9.58 8.24 10.22 ;
			RECT 7.6 2.78 8.24 10.22 ;
			RECT 1.82 1.98 2.46 3.26 ;

		END 

		ANTENNADIFFAREA 4.253 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 10.08 13.68 ;
			RECT 3.2 10.7 3.84 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 10.08 1.46 ;
			RECT 4.34 -0.48 6.56 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1.8 9.7 5.24 10.18 ;
			RECT 1.8 9.7 2.44 10.62 ;
			RECT 4.6 9.7 5.24 10.62 ;
			RECT 0.42 1.98 1.06 2.66 ;
			RECT 0.54 1.98 1.06 4.32 ;
			RECT 0.54 3.78 5.98 4.32 ;
			RECT 5.34 3.78 5.98 4.42 ;
			RECT 0.4 8.7 6.64 9.18 ;
			RECT 6 8.7 6.64 11.22 ;
			RECT 0.4 8.7 1.04 11.22 ;
			RECT 8.8 8.78 9.44 11.22 ;
			RECT 6 10.74 9.44 11.22 ;

	END

END AND222OXL

MACRO AND222O
	CLASS CORE ;
	FOREIGN AND222O 0 0  ;
	ORIGIN 0 0 ;
	SIZE 20.16 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 4.96 6.36 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.779 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 2.28 3.64 3.92 4.28 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.779 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 8.04 6.28 9.68 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.779 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 10.48 4.96 11.12 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.779 LAYER MTL1  ;
	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 13.36 3.96 14 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.779 LAYER MTL1  ;
	END E
	PIN F
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 11.92 6.28 12.56 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.779 LAYER MTL1  ;
	END F
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 17.2 7.54 17.94 10.18 ;
			RECT 14.46 7.54 17.94 8.02 ;
			RECT 14.8 2.08 15.44 8.02 ;
			RECT 14.46 6.28 15.1 10.18 ;
			RECT 9 2.9 15.44 3.38 ;
			RECT 13.8 2.08 15.44 3.38 ;
			RECT 9 2.12 9.64 3.38 ;

		END 

		ANTENNADIFFAREA 9.541 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 20.16 13.68 ;
			RECT 4.6 9.44 5.24 13.68 ;
			RECT 1.8 9.44 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 20.16 1.46 ;
			RECT 11.4 -0.48 12.04 2.36 ;
			RECT 6.58 -0.48 7.22 2.36 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 8.44 12.26 8.92 ;
			RECT 8.8 8.44 9.44 10.18 ;
			RECT 11.62 8.44 12.26 10.18 ;
			RECT 0.4 8.44 1.04 11.22 ;
			RECT 3.2 8.44 3.84 11.22 ;
			RECT 6 8.44 6.64 11.22 ;
			RECT 7.38 9.44 8.04 11.18 ;
			RECT 10.2 9.44 10.84 11.18 ;
			RECT 13.06 8.54 13.72 11.18 ;
			RECT 15.86 8.54 16.5 11.18 ;
			RECT 18.66 8.52 19.3 11.18 ;
			RECT 7.38 10.7 19.3 11.18 ;

	END

END AND222O

MACRO AND221OXL
	CLASS CORE ;
	FOREIGN AND221OXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 10.08 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.96 2.48 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.253 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.72 6.28 4.36 7.92 ;
			RECT 3.28 6.28 4.36 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.253 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 3.64 1.04 4.28 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.253 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 6.16 4.96 6.8 6.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.253 LAYER MTL1  ;
	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 9.04 7.6 9.68 9.26 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.181 LAYER MTL1  ;
	END E
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.4 9.56 8.24 11.22 ;
			RECT 7.6 3.28 8.24 11.22 ;
			RECT 1.94 3.78 8.24 4.26 ;
			RECT 7.58 3.28 8.24 4.26 ;
			RECT 1.94 2.98 2.58 4.26 ;

		END 

		ANTENNADIFFAREA 4.706 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 10.08 13.68 ;
			RECT 3.2 10.44 3.84 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 10.08 1.46 ;
			RECT 7.58 -0.48 8.22 2.26 ;
			RECT 4.58 -0.48 5.22 2.26 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 1.8 9.44 5.24 9.92 ;
			RECT 1.8 9.44 2.44 10.54 ;
			RECT 4.6 9.44 5.24 10.54 ;
			RECT 0.4 8.44 6.64 8.92 ;
			RECT 0.4 8.44 1.04 11.22 ;
			RECT 6 8.44 6.64 11.22 ;
			RECT 0.42 1.98 3.7 2.46 ;
			RECT 0.42 1.98 1.06 2.66 ;
			RECT 3.22 1.98 3.7 3.26 ;
			RECT 6.14 2.02 6.78 3.26 ;
			RECT 3.22 2.78 6.78 3.26 ;

	END

END AND221OXL

MACRO AND221O
	CLASS CORE ;
	FOREIGN AND221O 0 0  ;
	ORIGIN 0 0 ;
	SIZE 17.28 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 4.96 6.36 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.779 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 2.28 3.64 3.92 4.28 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.779 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 8.04 6.28 9.68 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.779 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 10.48 4.96 11.12 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.779 LAYER MTL1  ;
	END D
	PIN E
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 12.08 6.28 12.72 7.92 ;
			RECT 11.92 6.28 12.72 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.578 LAYER MTL1  ;
	END E
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 14.46 6.44 15.1 10.18 ;
			RECT 13.36 6.44 15.1 6.92 ;
			RECT 13.36 2.08 14 6.92 ;
			RECT 8.16 2.9 14 3.38 ;
			RECT 12 2.08 14 3.38 ;
			RECT 8.16 2.12 8.8 3.38 ;

		END 

		ANTENNADIFFAREA 5.874 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 17.28 13.68 ;
			RECT 4.6 9.44 5.24 13.68 ;
			RECT 1.8 9.44 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 17.28 1.46 ;
			RECT 10.56 -0.48 11.2 2.36 ;
			RECT 5.76 -0.48 6.4 2.36 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 8.44 12.26 8.92 ;
			RECT 8.8 8.44 9.44 10.18 ;
			RECT 11.62 8.44 12.26 10.18 ;
			RECT 0.4 8.44 1.04 11.22 ;
			RECT 3.2 8.44 3.84 11.22 ;
			RECT 6 8.44 6.64 11.22 ;
			RECT 7.38 9.44 8.04 11.18 ;
			RECT 10.2 9.44 10.84 11.18 ;
			RECT 13.06 8.54 13.72 11.18 ;
			RECT 15.82 8.54 16.5 11.18 ;
			RECT 7.38 10.7 16.5 11.18 ;

	END

END AND221O

MACRO AND22
	CLASS CORE ;
	FOREIGN AND22 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 7.54 1.04 9.18 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.08 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 5.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.08 LAYER MTL1  ;
	END B
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.64 8.94 5.36 11.22 ;
			RECT 4.72 1.98 5.36 11.22 ;
			RECT 4.24 1.98 5.36 3.62 ;

		END 

		ANTENNADIFFAREA 4.467 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 6.04 9.7 6.68 13.68 ;
			RECT 3.2 10.7 3.84 13.68 ;
			RECT 0.4 9.7 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 2.8 -0.48 3.44 2.62 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 1.98 1.04 3.62 ;
			RECT 0.4 3.14 3.72 3.62 ;
			RECT 3.24 3.14 3.72 5.78 ;
			RECT 3.64 4.14 4.12 10.18 ;
			RECT 1.8 9.7 4.12 10.18 ;
			RECT 1.8 9.7 2.44 10.9 ;

	END

END AND22

MACRO AND21OXL
	CLASS CORE ;
	FOREIGN AND21OXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 5.76 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 7.6 1.04 8.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.965 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 6.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.965 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 4.96 3.92 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.893 LAYER MTL1  ;
	END C
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.6 9.58 5.36 11.22 ;
			RECT 4.72 1.98 5.36 11.22 ;
			RECT 0.4 3.14 5.36 3.62 ;
			RECT 4.44 1.98 5.36 3.62 ;
			RECT 0.4 1.98 1.04 3.62 ;

		END 

		ANTENNADIFFAREA 3.022 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 5.76 13.68 ;
			RECT 1.8 10.7 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 5.76 1.46 ;
			RECT 2.8 -0.48 3.44 2.62 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 9.58 3.84 10.14 ;
			RECT 0.4 9.58 1.04 11.22 ;
			RECT 3.2 9.58 3.84 11.22 ;

	END

END AND21OXL

MACRO AND21O
	CLASS CORE ;
	FOREIGN AND21O 0 0  ;
	ORIGIN 0 0 ;
	SIZE 8.64 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 3.96 1.04 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.261 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 2.28 6.28 3.92 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.261 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 4.96 5.64 5.6 ;
			RECT 5 3.96 5.64 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.059 LAYER MTL1  ;
	END C
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 5.54 10.58 7.48 11.22 ;
			RECT 6.16 2.96 6.8 11.22 ;
			RECT 4 2.96 6.8 3.44 ;
			RECT 4 1.98 4.88 3.44 ;
			RECT 1.68 3.14 4.48 3.62 ;
			RECT 0.4 2.96 2.16 3.44 ;
			RECT 0.4 2.34 1.04 3.44 ;

		END 

		ANTENNADIFFAREA 6.48 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 8.64 13.68 ;
			RECT 3.12 9.76 3.76 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 8.64 1.46 ;
			RECT 2.8 -0.48 3.44 2.62 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 2.12 8.76 5.18 9.24 ;
			RECT 4.54 8.76 5.18 9.8 ;
			RECT 2.12 8.76 2.6 11.22 ;
			RECT 0.4 10.58 2.6 11.22 ;

	END

END AND21O

MACRO AND211OXL
	CLASS CORE ;
	FOREIGN AND211OXL 0 0  ;
	ORIGIN 0 0 ;
	SIZE 7.2 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 4.96 2.48 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.253 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 3.64 1.04 4.28 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.253 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 6.28 3.92 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.181 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.72 3.98 5.36 5.62 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 1.181 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 5.6 8.76 6.8 11.22 ;
			RECT 6.16 1.98 6.8 11.22 ;
			RECT 2.82 2.78 6.8 3.26 ;
			RECT 6.1 1.98 6.8 3.26 ;
			RECT 2.82 1.98 3.46 3.26 ;

		END 

		ANTENNADIFFAREA 3.872 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 7.2 13.68 ;
			RECT 1.8 9.76 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 7.2 1.46 ;
			RECT 4.46 -0.48 5.1 2.26 ;
			RECT 0.42 -0.48 1.06 2.62 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 8.76 3.84 9.24 ;
			RECT 0.4 8.76 1.04 11.22 ;
			RECT 3.2 8.76 3.84 11.22 ;

	END

END AND211OXL

MACRO AND211O
	CLASS CORE ;
	FOREIGN AND211O 0 0  ;
	ORIGIN 0 0 ;
	SIZE 14.4 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 3.28 4.96 4.92 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.779 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.84 3.64 2.48 4.28 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.779 LAYER MTL1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 7.6 6.28 9.24 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.578 LAYER MTL1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 10.48 3.96 11.12 5.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 2.578 LAYER MTL1  ;
	END D
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 11.92 2.12 12.56 9.56 ;
			RECT 11.64 8.58 12.28 10.22 ;
			RECT 8.08 2.9 12.56 3.38 ;
			RECT 11 2.12 12.56 3.38 ;
			RECT 8.08 2.12 8.72 3.38 ;

		END 

		ANTENNADIFFAREA 5.918 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 14.4 13.68 ;
			RECT 4.6 9.44 5.24 13.68 ;
			RECT 1.8 9.44 2.44 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 14.4 1.46 ;
			RECT 9.6 -0.48 10.24 2.36 ;
			RECT 5.68 -0.48 6.32 2.86 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 8.44 9.48 8.92 ;
			RECT 8.84 8.44 9.48 10.22 ;
			RECT 0.4 8.44 1.04 11.22 ;
			RECT 3.2 8.44 3.84 11.22 ;
			RECT 6 8.44 6.64 11.22 ;
			RECT 7.44 9.44 8.08 11.22 ;
			RECT 10.24 8.44 10.88 11.22 ;
			RECT 13.08 8.44 13.72 11.22 ;
			RECT 7.44 10.74 13.72 11.22 ;

	END

END AND211O

MACRO AND2
	CLASS CORE ;
	FOREIGN AND2 0 0  ;
	ORIGIN 0 0 ;
	SIZE 5.76 BY 13.2 ;
	SYMMETRY X Y ;
	SITE standard ;
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 0.4 7.6 1.04 9.24 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.72 LAYER MTL1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 1.84 5.28 2.48 6.92 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAGATEAREA 0.72 LAYER MTL1  ;
	END B
	PIN O
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER MTL1 ;
			RECT 4.64 8.94 5.36 11.22 ;
			RECT 4.72 1.98 5.36 11.22 ;
			RECT 4.24 1.98 5.36 2.62 ;

		END 

		ANTENNADIFFAREA 3.098 LAYER MTL1  ;
	END O
	PIN vddd!
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 11.74 5.76 13.68 ;
			RECT 3.2 10.22 3.84 13.68 ;
			RECT 0.4 10.22 1.04 13.68 ;

		END 

	END vddd!
	PIN gndd!
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER MTL1 ;
			RECT 0 -0.48 5.76 1.46 ;
			RECT 2.8 -0.48 3.44 2.62 ;

		END 

	END gndd!
	OBS
			LAYER MTL1 ;
			RECT 0.4 1.98 1.04 3.62 ;
			RECT 0.4 3.14 4.12 3.62 ;
			RECT 3.48 3.14 4.12 5.02 ;
			RECT 3.56 3.14 4.12 9.7 ;
			RECT 1.8 9.22 4.12 9.7 ;
			RECT 1.8 9.22 2.44 11.22 ;

	END

END AND2

END LIBRARY
