// 
//	raifes_gpio
//
`include "raifes_hasti_constants.vh"

`define GPIO_BASE_ADDR	32'hC0000000

module raifes_gpio(
		// system clk and reset
		input			reset,
		input			clk,

		// gpio in/outputs
		output	reg	[7:0]	gpio_d,
		output	reg	[7:0]	gpio_en,
		input		[7:0]	gpio_i,

		// system bus 
	        input	[`HASTI_ADDR_WIDTH-1:0]  haddr,
        	input				hwrite,			// unused, as imem is read-only (typically)
	        input	[`HASTI_SIZE_WIDTH-1:0]  hsize,
		input	[`HASTI_BURST_WIDTH-1:0] hburst,
	        input 			   	hmastlock,
	        input	[`HASTI_PROT_WIDTH-1:0]  hprot,
	        input	[`HASTI_TRANS_WIDTH-1:0] htrans,
	        input	[`HASTI_BUS_WIDTH-1:0]   hwdata,			// unused, as imem is read-only (typically)
	        output	reg	[`HASTI_BUS_WIDTH-1:0]    hrdata,
	        output 	reg			   	hready,
	        output	reg	[`HASTI_RESP_WIDTH-1:0]   hresp
);


`define GPIO_IDLE 0
`define GPIO_READ_D 1
`define GPIO_READ_EN 2
`define GPIO_WRITE_D 3
`define GPIO_WRITE_EN 4

reg	[2:0]	state, next_state;
reg	[`HASTI_ADDR_WIDTH-1:0]	addr_r;	// hold addr in case of write operations

always @(posedge clk) begin
	if(reset) begin 
		state <= `GPIO_IDLE;
	end else begin
		state <= next_state;


		if(next_state == `GPIO_READ_D) begin
			hrdata <= {gpio_i,gpio_i,gpio_i,gpio_i};
		end else
		if(next_state == `GPIO_READ_EN) begin
			hrdata <= {gpio_en,gpio_en,gpio_en,gpio_en};
		end else
		if(state == `GPIO_WRITE_D) begin
			gpio_d <= hwdata[7:0];
		end else
		if(state == `GPIO_WRITE_EN) begin
			gpio_en <= hwdata[7:0];
		end
	end
end

always @(*) begin
	hready = 1'b0;
	case (state) 
		`GPIO_IDLE	:	begin
					hready = 1'b1;
					if((haddr == `GPIO_BASE_ADDR) && |htrans) begin
						next_state = |hwrite ? `GPIO_WRITE_D : `GPIO_READ_D;
					end else 
					if((haddr == `GPIO_BASE_ADDR+4) && |htrans) begin
						next_state = |hwrite ? `GPIO_WRITE_EN : `GPIO_READ_EN;
					end else next_state = `GPIO_IDLE;
				end
		`GPIO_READ_D	:	begin
					next_state = `GPIO_IDLE;		
				end
		`GPIO_WRITE_D :	begin
					next_state = `GPIO_IDLE;
				end
		`GPIO_READ_EN : 	begin 
					next_state = `GPIO_IDLE;
				end
		`GPIO_WRITE_EN :	begin 
					next_state = `GPIO_IDLE;
				end
	endcase
end

endmodule
